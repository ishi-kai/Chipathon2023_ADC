* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt TOP VDD Vctrl GND Vin Vout
X0 Vout.t18 a_n2515_0.t10 Vin.t5 VDD.t21 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1 a_n2515_0.t4 Vctrl.t0 GND.t29 GND.t28 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2 a_n2515_0.t5 Vctrl.t1 GND.t27 GND.t26 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3 VDD.t3 Vctrl.t2 a_n2515_0.t1 VDD.t2 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4 Vin.t8 a_n2515_0.t11 Vout.t17 VDD.t20 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X5 Vin.t11 a_n2515_0.t12 Vout.t16 VDD.t19 pfet_03v3 ad=1.82p pd=6.9u as=0.728p ps=3.32u w=2.8u l=0.28u
X6 GND.t25 Vctrl.t3 a_n2515_0.t5 GND.t24 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X7 Vout.t6 a_n2515_0.t13 GND.t49 GND.t48 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X8 Vout.t19 a_n2515_0.t14 GND.t47 GND.t46 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X9 Vout.t15 a_n2515_0.t15 Vin.t3 VDD.t18 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X10 GND.t45 a_n2515_0.t16 Vout.t22 GND.t44 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X11 VDD.t5 Vctrl.t4 a_n2515_0.t3 VDD.t4 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X12 Vout.t21 a_n2515_0.t17 GND.t43 GND.t42 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X13 a_n2515_0.t1 Vctrl.t5 VDD.t7 VDD.t6 pfet_03v3 ad=0.728p pd=3.32u as=1.82p ps=6.9u w=2.8u l=0.28u
X14 a_n2515_0.t0 Vctrl.t6 VDD.t9 VDD.t8 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X15 VDD.t23 Vctrl.t7 a_n2515_0.t8 VDD.t22 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X16 Vout.t14 a_n2515_0.t18 Vin.t6 VDD.t17 pfet_03v3 ad=0.728p pd=3.32u as=1.82p ps=6.9u w=2.8u l=0.28u
X17 Vout.t13 a_n2515_0.t19 Vin.t7 VDD.t16 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X18 Vin.t9 a_n2515_0.t20 Vout.t12 VDD.t15 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X19 Vout.t29 Vctrl.t8 Vin.t19 GND.t23 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X20 a_n2515_0.t9 Vctrl.t9 GND.t22 GND.t21 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X21 Vin.t16 Vctrl.t10 Vout.t26 GND.t20 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X22 Vin.t15 Vctrl.t11 Vout.t25 GND.t19 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X23 GND.t18 Vctrl.t12 a_n2515_0.t9 GND.t17 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X24 GND.t16 Vctrl.t13 a_n2515_0.t6 GND.t15 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X25 Vin.t14 Vctrl.t14 Vout.t24 GND.t14 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X26 a_n2515_0.t2 Vctrl.t15 GND.t13 GND.t12 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X27 Vout.t27 Vctrl.t16 Vin.t17 GND.t11 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X28 GND.t10 Vctrl.t17 a_n2515_0.t4 GND.t9 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X29 GND.t41 a_n2515_0.t21 Vout.t3 GND.t40 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X30 Vout.t7 a_n2515_0.t22 GND.t39 GND.t38 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X31 a_n2515_0.t3 Vctrl.t18 VDD.t27 VDD.t26 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X32 GND.t37 a_n2515_0.t23 Vout.t4 GND.t36 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X33 Vin.t10 a_n2515_0.t24 Vout.t11 VDD.t14 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X34 a_n2515_0.t8 Vctrl.t19 VDD.t25 VDD.t24 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X35 VDD.t29 Vctrl.t20 a_n2515_0.t7 VDD.t28 pfet_03v3 ad=1.82p pd=6.9u as=0.728p ps=3.32u w=2.8u l=0.28u
X36 GND.t35 a_n2515_0.t25 Vout.t8 GND.t34 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X37 Vout.t10 a_n2515_0.t26 Vin.t12 VDD.t13 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X38 Vout.t20 a_n2515_0.t27 GND.t33 GND.t32 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X39 Vin.t4 a_n2515_0.t28 Vout.t9 VDD.t12 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X40 Vout.t23 Vctrl.t21 Vin.t13 GND.t8 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X41 a_n2515_0.t7 Vctrl.t22 VDD.t11 VDD.t10 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X42 Vin.t0 Vctrl.t23 Vout.t0 GND.t7 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X43 VDD.t1 Vctrl.t24 a_n2515_0.t0 VDD.t0 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X44 Vout.t1 Vctrl.t25 Vin.t1 GND.t6 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X45 Vout.t2 Vctrl.t26 Vin.t2 GND.t5 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X46 a_n2515_0.t6 Vctrl.t27 GND.t4 GND.t3 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X47 GND.t2 Vctrl.t28 a_n2515_0.t2 GND.t1 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X48 Vin.t18 Vctrl.t29 Vout.t28 GND.t0 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X49 GND.t31 a_n2515_0.t29 Vout.t5 GND.t30 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
R0 a_n2515_0.n3 a_n2515_0.t18 56.0276
R1 a_n2515_0.n4 a_n2515_0.t29 56.019
R2 a_n2515_0.n3 a_n2515_0.t24 55.9719
R3 a_n2515_0.n3 a_n2515_0.t19 55.9719
R4 a_n2515_0.n3 a_n2515_0.t11 55.9719
R5 a_n2515_0.n3 a_n2515_0.t10 55.9719
R6 a_n2515_0.n3 a_n2515_0.t28 55.9719
R7 a_n2515_0.n0 a_n2515_0.t26 55.9719
R8 a_n2515_0.n0 a_n2515_0.t20 55.9719
R9 a_n2515_0.n0 a_n2515_0.t15 55.9719
R10 a_n2515_0.n0 a_n2515_0.t12 55.9719
R11 a_n2515_0.n4 a_n2515_0.t27 55.9719
R12 a_n2515_0.n4 a_n2515_0.t25 55.9719
R13 a_n2515_0.n4 a_n2515_0.t17 55.9719
R14 a_n2515_0.n4 a_n2515_0.t23 55.9719
R15 a_n2515_0.n4 a_n2515_0.t22 55.9719
R16 a_n2515_0.n4 a_n2515_0.t16 55.9719
R17 a_n2515_0.n4 a_n2515_0.t13 55.9719
R18 a_n2515_0.n4 a_n2515_0.t21 55.9719
R19 a_n2515_0.n4 a_n2515_0.t14 55.9719
R20 a_n2515_0.n1 a_n2515_0.t9 3.87048
R21 a_n2515_0.n1 a_n2515_0.t6 3.68704
R22 a_n2515_0.n1 a_n2515_0.t2 3.68704
R23 a_n2515_0.n1 a_n2515_0.t4 3.68704
R24 a_n2515_0.n1 a_n2515_0.t5 3.68704
R25 a_n2515_0.n2 a_n2515_0.t1 3.53719
R26 a_n2515_0.n2 a_n2515_0.t7 3.37808
R27 a_n2515_0.n2 a_n2515_0.t8 3.37808
R28 a_n2515_0.n2 a_n2515_0.t3 3.37808
R29 a_n2515_0.t0 a_n2515_0.n2 3.37783
R30 a_n2515_0.n2 a_n2515_0.n1 1.83641
R31 a_n2515_0.n0 a_n2515_0.n4 1.82216
R32 a_n2515_0.n2 a_n2515_0.n0 1.29508
R33 a_n2515_0.n0 a_n2515_0.n3 1.12477
R34 Vin.n0 Vin.t14 15.8618
R35 Vin.n9 Vin.t1 15.8393
R36 Vin.n0 Vin.t11 15.7537
R37 Vin.n9 Vin.t6 15.7496
R38 Vin.n11 Vin.n10 14.963
R39 Vin.n15 Vin.n14 14.9583
R40 Vin.n4 Vin.n3 14.9559
R41 Vin.n6 Vin.n5 14.9547
R42 Vin.n13 Vin.n12 14.7096
R43 Vin.n17 Vin.n16 14.7035
R44 Vin.n8 Vin.n7 14.7035
R45 Vin.n2 Vin.n1 14.6941
R46 Vin.n12 Vin.t7 0.6505
R47 Vin.n12 Vin.t10 0.6505
R48 Vin.n16 Vin.t5 0.6505
R49 Vin.n16 Vin.t8 0.6505
R50 Vin.n7 Vin.t12 0.6505
R51 Vin.n7 Vin.t4 0.6505
R52 Vin.n1 Vin.t3 0.6505
R53 Vin.n1 Vin.t9 0.6505
R54 Vin.n10 Vin.t2 0.5855
R55 Vin.n10 Vin.t16 0.5855
R56 Vin.n14 Vin.t19 0.5855
R57 Vin.n14 Vin.t15 0.5855
R58 Vin.n5 Vin.t13 0.5855
R59 Vin.n5 Vin.t0 0.5855
R60 Vin.n3 Vin.t17 0.5855
R61 Vin.n3 Vin.t18 0.5855
R62 Vin.n11 Vin.n9 0.0340106
R63 Vin.n2 Vin.n0 0.0332447
R64 Vin.n6 Vin.n4 0.031234
R65 Vin.n15 Vin.n13 0.0308511
R66 Vin Vin.n8 0.0243404
R67 Vin Vin.n17 0.00653191
R68 Vin.n4 Vin.n2 0.000978723
R69 Vin.n17 Vin.n15 0.000882979
R70 Vin.n8 Vin.n6 0.000691489
R71 Vin.n13 Vin.n11 0.000595745
R72 Vout.n21 Vout.n19 10.5979
R73 Vout.n12 Vout.n10 10.553
R74 Vout.n21 Vout.n20 10.4369
R75 Vout.n27 Vout.n26 10.4308
R76 Vout.n25 Vout.n24 10.4308
R77 Vout.n23 Vout.n22 10.4308
R78 Vout.n12 Vout.n11 10.4156
R79 Vout.n16 Vout.n15 10.4129
R80 Vout.n14 Vout.n13 10.4121
R81 Vout.n18 Vout.n17 10.4121
R82 Vout.n2 Vout.n0 10.357
R83 Vout.n4 Vout.n3 10.2004
R84 Vout.n8 Vout.n7 10.2004
R85 Vout.n6 Vout.n5 10.198
R86 Vout.n2 Vout.n1 10.1921
R87 Vout.n28 Vout.n9 2.3885
R88 Vout.n0 Vout.t11 0.6505
R89 Vout.n0 Vout.t14 0.6505
R90 Vout.n1 Vout.t17 0.6505
R91 Vout.n1 Vout.t13 0.6505
R92 Vout.n3 Vout.t9 0.6505
R93 Vout.n3 Vout.t18 0.6505
R94 Vout.n5 Vout.t12 0.6505
R95 Vout.n5 Vout.t10 0.6505
R96 Vout.n7 Vout.t16 0.6505
R97 Vout.n7 Vout.t15 0.6505
R98 Vout.n10 Vout.t26 0.5855
R99 Vout.n10 Vout.t1 0.5855
R100 Vout.n11 Vout.t25 0.5855
R101 Vout.n11 Vout.t2 0.5855
R102 Vout.n13 Vout.t0 0.5855
R103 Vout.n13 Vout.t29 0.5855
R104 Vout.n15 Vout.t28 0.5855
R105 Vout.n15 Vout.t23 0.5855
R106 Vout.n17 Vout.t24 0.5855
R107 Vout.n17 Vout.t27 0.5855
R108 Vout.n26 Vout.t8 0.5855
R109 Vout.n26 Vout.t20 0.5855
R110 Vout.n24 Vout.t4 0.5855
R111 Vout.n24 Vout.t21 0.5855
R112 Vout.n22 Vout.t22 0.5855
R113 Vout.n22 Vout.t7 0.5855
R114 Vout.n20 Vout.t3 0.5855
R115 Vout.n20 Vout.t6 0.5855
R116 Vout.n19 Vout.t5 0.5855
R117 Vout.n19 Vout.t19 0.5855
R118 Vout.n9 Vout.n8 0.528502
R119 Vout.n29 Vout.n18 0.364991
R120 Vout.n28 Vout.n27 0.2945
R121 Vout Vout.n29 0.263973
R122 Vout.n8 Vout.n6 0.161
R123 Vout.n6 Vout.n4 0.1605
R124 Vout.n4 Vout.n2 0.1605
R125 Vout.n25 Vout.n23 0.1605
R126 Vout.n27 Vout.n25 0.1605
R127 Vout.n23 Vout.n21 0.1585
R128 Vout.n18 Vout.n16 0.139126
R129 Vout.n14 Vout.n12 0.136566
R130 Vout.n16 Vout.n14 0.13486
R131 Vout Vout.n9 0.00767791
R132 Vout.n29 Vout.n28 0.00376492
R133 VDD VDD.t19 312.592
R134 VDD.n0 VDD.t28 311.132
R135 VDD.t28 VDD.t10 191.388
R136 VDD.t10 VDD.t22 191.388
R137 VDD.t22 VDD.t24 191.388
R138 VDD.t24 VDD.t0 191.388
R139 VDD.t0 VDD.t8 191.388
R140 VDD.t8 VDD.t4 191.388
R141 VDD.t4 VDD.t26 191.388
R142 VDD.t26 VDD.t2 191.388
R143 VDD.t2 VDD.t6 191.388
R144 VDD.t19 VDD.t18 191.388
R145 VDD.t18 VDD.t15 191.388
R146 VDD.t15 VDD.t13 191.388
R147 VDD.t13 VDD.t12 191.388
R148 VDD.t12 VDD.t21 191.388
R149 VDD.t21 VDD.t20 191.388
R150 VDD.t20 VDD.t16 191.388
R151 VDD.t16 VDD.t14 191.388
R152 VDD.t14 VDD.t17 191.388
R153 VDD.n5 VDD.t7 2.95135
R154 VDD.n0 VDD.t29 2.0905
R155 VDD.n5 VDD.n4 1.80644
R156 VDD.n6 VDD.n3 1.80644
R157 VDD.n7 VDD.n2 1.80644
R158 VDD.n8 VDD.n1 1.80644
R159 VDD.n4 VDD.t27 0.6505
R160 VDD.n4 VDD.t3 0.6505
R161 VDD.n3 VDD.t9 0.6505
R162 VDD.n3 VDD.t5 0.6505
R163 VDD.n2 VDD.t25 0.6505
R164 VDD.n2 VDD.t1 0.6505
R165 VDD.n1 VDD.t11 0.6505
R166 VDD.n1 VDD.t23 0.6505
R167 VDD.n9 VDD.n0 0.261581
R168 VDD VDD.n9 0.145415
R169 VDD.n9 VDD.n8 0.131992
R170 VDD.n8 VDD.n7 0.0981271
R171 VDD.n7 VDD.n6 0.0981271
R172 VDD.n6 VDD.n5 0.0981271
R173 Vctrl.n10 Vctrl.t20 56.1018
R174 Vctrl.n0 Vctrl.t14 56.0719
R175 Vctrl.n9 Vctrl.t3 56.0141
R176 Vctrl.n15 Vctrl.t5 55.9719
R177 Vctrl.n16 Vctrl.t2 55.9719
R178 Vctrl.n17 Vctrl.t18 55.9719
R179 Vctrl.n18 Vctrl.t4 55.9719
R180 Vctrl.n19 Vctrl.t6 55.9719
R181 Vctrl.n14 Vctrl.t24 55.9719
R182 Vctrl.n13 Vctrl.t19 55.9719
R183 Vctrl.n12 Vctrl.t7 55.9719
R184 Vctrl.n11 Vctrl.t22 55.9719
R185 Vctrl.n15 Vctrl.t9 55.9719
R186 Vctrl.n16 Vctrl.t12 55.9719
R187 Vctrl.n17 Vctrl.t27 55.9719
R188 Vctrl.n18 Vctrl.t13 55.9719
R189 Vctrl.n19 Vctrl.t15 55.9719
R190 Vctrl.n14 Vctrl.t28 55.9719
R191 Vctrl.n13 Vctrl.t0 55.9719
R192 Vctrl.n12 Vctrl.t17 55.9719
R193 Vctrl.n11 Vctrl.t1 55.9719
R194 Vctrl.n8 Vctrl.t25 55.9719
R195 Vctrl.n7 Vctrl.t10 55.9719
R196 Vctrl.n6 Vctrl.t26 55.9719
R197 Vctrl.n5 Vctrl.t11 55.9719
R198 Vctrl.n4 Vctrl.t8 55.9719
R199 Vctrl.n3 Vctrl.t23 55.9719
R200 Vctrl.n2 Vctrl.t21 55.9719
R201 Vctrl.n1 Vctrl.t29 55.9719
R202 Vctrl.n0 Vctrl.t16 55.9719
R203 Vctrl.n9 Vctrl.n8 0.7055
R204 Vctrl.n1 Vctrl.n0 0.1005
R205 Vctrl.n2 Vctrl.n1 0.1005
R206 Vctrl.n3 Vctrl.n2 0.1005
R207 Vctrl.n4 Vctrl.n3 0.1005
R208 Vctrl.n5 Vctrl.n4 0.1005
R209 Vctrl.n6 Vctrl.n5 0.1005
R210 Vctrl.n7 Vctrl.n6 0.1005
R211 Vctrl.n8 Vctrl.n7 0.1005
R212 Vctrl.n10 Vctrl.n9 0.0961962
R213 Vctrl.n12 Vctrl.n11 0.0475588
R214 Vctrl.n13 Vctrl.n12 0.0475588
R215 Vctrl.n14 Vctrl.n13 0.0475588
R216 Vctrl.n19 Vctrl.n18 0.0475588
R217 Vctrl.n18 Vctrl.n17 0.0475588
R218 Vctrl.n17 Vctrl.n16 0.0475588
R219 Vctrl.n16 Vctrl.n15 0.0475588
R220 Vctrl.n11 Vctrl.n10 0.0363824
R221 Vctrl Vctrl.n14 0.0334412
R222 Vctrl Vctrl.n19 0.0146176
R223 GND.t21 GND.n17 24415
R224 GND.n17 GND.n16 14963.3
R225 GND.n17 GND.n4 6221
R226 GND.t6 GND.n4 1245.51
R227 GND.n18 GND.n4 993.961
R228 GND.n16 GND.t32 867.15
R229 GND.n18 GND.t24 613.208
R230 GND.n15 GND.t14 608.159
R231 GND.n16 GND.n15 467.067
R232 GND.t24 GND.t26 392.454
R233 GND.t26 GND.t9 392.454
R234 GND.t9 GND.t28 392.454
R235 GND.t28 GND.t1 392.454
R236 GND.t1 GND.t12 392.454
R237 GND.t12 GND.t15 392.454
R238 GND.t15 GND.t3 392.454
R239 GND.t3 GND.t17 392.454
R240 GND.t17 GND.t21 392.454
R241 GND.t14 GND.t11 389.223
R242 GND.t11 GND.t0 389.223
R243 GND.t0 GND.t8 389.223
R244 GND.t8 GND.t7 389.223
R245 GND.t7 GND.t23 389.223
R246 GND.t23 GND.t19 389.223
R247 GND.t19 GND.t5 389.223
R248 GND.t5 GND.t20 389.223
R249 GND.t20 GND.t6 389.223
R250 GND.t30 GND.n14 308.666
R251 GND.t46 GND.t30 193.238
R252 GND.t40 GND.t46 193.238
R253 GND.t48 GND.t40 193.238
R254 GND.t44 GND.t48 193.238
R255 GND.t38 GND.t44 193.238
R256 GND.t36 GND.t38 193.238
R257 GND.t42 GND.t36 193.238
R258 GND.t34 GND.t42 193.238
R259 GND.t32 GND.t34 193.238
R260 GND.n9 GND.t33 7.21552
R261 GND.n14 GND.t31 6.80897
R262 GND.n12 GND.n6 6.31687
R263 GND.n11 GND.n7 6.31687
R264 GND.n13 GND.n5 6.3142
R265 GND.n10 GND.n8 6.31016
R266 GND.n24 GND.n23 4.61975
R267 GND.n20 GND.n1 4.61975
R268 GND.n21 GND.n20 4.5005
R269 GND.n23 GND.n22 4.5005
R270 GND.n29 GND.t22 3.91509
R271 GND.n15 GND.n0 3.68746
R272 GND.n32 GND.n25 2.90641
R273 GND.n31 GND.n26 2.90641
R274 GND.n30 GND.n27 2.90641
R275 GND.n29 GND.n28 2.90641
R276 GND.n19 GND.n3 2.33691
R277 GND.n3 GND.n2 2.33309
R278 GND.n2 GND.t25 2.1605
R279 GND.n19 GND.n18 2.0805
R280 GND GND.n0 0.703625
R281 GND.n5 GND.t47 0.5855
R282 GND.n5 GND.t41 0.5855
R283 GND.n6 GND.t49 0.5855
R284 GND.n6 GND.t45 0.5855
R285 GND.n7 GND.t39 0.5855
R286 GND.n7 GND.t37 0.5855
R287 GND.n8 GND.t43 0.5855
R288 GND.n8 GND.t35 0.5855
R289 GND.n25 GND.t27 0.5855
R290 GND.n25 GND.t10 0.5855
R291 GND.n26 GND.t29 0.5855
R292 GND.n26 GND.t2 0.5855
R293 GND.n27 GND.t13 0.5855
R294 GND.n27 GND.t16 0.5855
R295 GND.n28 GND.t4 0.5855
R296 GND.n28 GND.t18 0.5855
R297 GND.n14 GND.n13 0.28617
R298 GND.n9 GND.n0 0.263882
R299 GND.n33 GND.n24 0.220767
R300 GND GND.n33 0.185132
R301 GND.n33 GND.n32 0.139801
R302 GND.n10 GND.n9 0.115978
R303 GND.n11 GND.n10 0.106382
R304 GND.n30 GND.n29 0.106382
R305 GND.n13 GND.n12 0.106051
R306 GND.n32 GND.n31 0.106051
R307 GND.n12 GND.n11 0.105721
R308 GND.n31 GND.n30 0.105721
R309 GND.n23 GND.n2 0.066875
R310 GND.n20 GND.n19 0.064625
R311 GND.n21 GND.n3 0.0539756
R312 GND.n22 GND.n1 0.0426622
R313 GND.n22 GND.n21 0.00131081
R314 GND.n24 GND.n1 0.00131081
C0 Vin VDD 0.64647f
C1 Vctrl VDD 1.73327f
C2 Vout Vin 7.27658f
C3 Vout Vctrl 0.576084f
C4 Vctrl Vin 0.85985f
C5 Vout VDD 0.33441f
C6 Vout GND 6.420404f
C7 Vin GND 2.003741f
C8 Vctrl GND 5.275005f
C9 VDD GND 17.525967f
C10 Vctrl.t20 GND 0.039242f
C11 Vctrl.t14 GND 0.039161f
C12 Vctrl.t16 GND 0.039019f
C13 Vctrl.n0 GND 0.134377f
C14 Vctrl.t29 GND 0.039019f
C15 Vctrl.n1 GND 0.054949f
C16 Vctrl.t21 GND 0.039019f
C17 Vctrl.n2 GND 0.054949f
C18 Vctrl.t23 GND 0.039019f
C19 Vctrl.n3 GND 0.054949f
C20 Vctrl.t8 GND 0.039019f
C21 Vctrl.n4 GND 0.054949f
C22 Vctrl.t11 GND 0.039019f
C23 Vctrl.n5 GND 0.054949f
C24 Vctrl.t26 GND 0.039019f
C25 Vctrl.n6 GND 0.054949f
C26 Vctrl.t10 GND 0.039019f
C27 Vctrl.n7 GND 0.054949f
C28 Vctrl.t25 GND 0.039019f
C29 Vctrl.n8 GND 0.165287f
C30 Vctrl.t3 GND 0.039038f
C31 Vctrl.n9 GND 0.161285f
C32 Vctrl.n10 GND 0.073488f
C33 Vctrl.t1 GND 0.039019f
C34 Vctrl.t22 GND 0.039169f
C35 Vctrl.n11 GND 0.106041f
C36 Vctrl.t17 GND 0.039019f
C37 Vctrl.t7 GND 0.039169f
C38 Vctrl.n12 GND 0.115245f
C39 Vctrl.t0 GND 0.039019f
C40 Vctrl.t19 GND 0.039169f
C41 Vctrl.n13 GND 0.115245f
C42 Vctrl.t28 GND 0.039019f
C43 Vctrl.t24 GND 0.039169f
C44 Vctrl.n14 GND 0.103619f
C45 Vctrl.t15 GND 0.039019f
C46 Vctrl.t13 GND 0.039019f
C47 Vctrl.t27 GND 0.039019f
C48 Vctrl.t12 GND 0.039019f
C49 Vctrl.t9 GND 0.039019f
C50 Vctrl.t5 GND 0.039169f
C51 Vctrl.n15 GND 0.095849f
C52 Vctrl.t2 GND 0.039169f
C53 Vctrl.n16 GND 0.115245f
C54 Vctrl.t18 GND 0.039169f
C55 Vctrl.n17 GND 0.115245f
C56 Vctrl.t4 GND 0.039169f
C57 Vctrl.n18 GND 0.115245f
C58 Vctrl.t6 GND 0.039169f
C59 Vctrl.n19 GND 0.088117f
C60 VDD.t17 GND 0.29116f
C61 VDD.t14 GND 0.123898f
C62 VDD.t16 GND 0.123898f
C63 VDD.t20 GND 0.123898f
C64 VDD.t21 GND 0.123898f
C65 VDD.t12 GND 0.123898f
C66 VDD.t13 GND 0.123898f
C67 VDD.t15 GND 0.123898f
C68 VDD.t18 GND 0.123898f
C69 VDD.t19 GND 0.165356f
C70 VDD.t6 GND 0.29116f
C71 VDD.t2 GND 0.123898f
C72 VDD.t26 GND 0.123898f
C73 VDD.t4 GND 0.123898f
C74 VDD.t8 GND 0.123898f
C75 VDD.t0 GND 0.123898f
C76 VDD.t24 GND 0.123898f
C77 VDD.t22 GND 0.123898f
C78 VDD.t10 GND 0.123898f
C79 VDD.t28 GND 0.163498f
C80 VDD.t29 GND 0.0445f
C81 VDD.n0 GND 0.307098f
C82 VDD.t11 GND 0.013486f
C83 VDD.t23 GND 0.013486f
C84 VDD.n1 GND 0.044291f
C85 VDD.t25 GND 0.013486f
C86 VDD.t1 GND 0.013486f
C87 VDD.n2 GND 0.044291f
C88 VDD.t9 GND 0.013486f
C89 VDD.t5 GND 0.013486f
C90 VDD.n3 GND 0.044291f
C91 VDD.t27 GND 0.013486f
C92 VDD.t3 GND 0.013486f
C93 VDD.n4 GND 0.044291f
C94 VDD.t7 GND 0.050177f
C95 VDD.n5 GND -0.177183f
C96 VDD.n6 GND 0.133881f
C97 VDD.n7 GND 0.133881f
C98 VDD.n8 GND 0.149046f
C99 VDD.n9 GND 0.191439f
C100 Vout.t11 GND 0.032704f
C101 Vout.t14 GND 0.032704f
C102 Vout.n0 GND 0.159978f
C103 Vout.t17 GND 0.032704f
C104 Vout.t13 GND 0.032704f
C105 Vout.n1 GND 0.1539f
C106 Vout.n2 GND 0.448318f
C107 Vout.t9 GND 0.032704f
C108 Vout.t18 GND 0.032704f
C109 Vout.n3 GND 0.155988f
C110 Vout.n4 GND 0.154881f
C111 Vout.t12 GND 0.032704f
C112 Vout.t10 GND 0.032704f
C113 Vout.n5 GND 0.155392f
C114 Vout.n6 GND 0.154997f
C115 Vout.t16 GND 0.032704f
C116 Vout.t15 GND 0.032704f
C117 Vout.n7 GND 0.155988f
C118 Vout.n8 GND 0.317081f
C119 Vout.n9 GND 0.242085f
C120 Vout.t26 GND 0.032704f
C121 Vout.t1 GND 0.032704f
C122 Vout.n10 GND 0.157478f
C123 Vout.t25 GND 0.032704f
C124 Vout.t2 GND 0.032704f
C125 Vout.n11 GND 0.152907f
C126 Vout.n12 GND 0.529333f
C127 Vout.t0 GND 0.032704f
C128 Vout.t29 GND 0.032704f
C129 Vout.n13 GND 0.15203f
C130 Vout.n14 GND 0.180901f
C131 Vout.t28 GND 0.032704f
C132 Vout.t23 GND 0.032704f
C133 Vout.n15 GND 0.153694f
C134 Vout.n16 GND 0.182582f
C135 Vout.t24 GND 0.032704f
C136 Vout.t27 GND 0.032704f
C137 Vout.n17 GND 0.15203f
C138 Vout.n18 GND 0.31784f
C139 Vout.t5 GND 0.032704f
C140 Vout.t19 GND 0.032704f
C141 Vout.n19 GND 0.160478f
C142 Vout.t3 GND 0.032704f
C143 Vout.t6 GND 0.032704f
C144 Vout.n20 GND 0.156394f
C145 Vout.n21 GND 0.421514f
C146 Vout.t22 GND 0.032704f
C147 Vout.t7 GND 0.032704f
C148 Vout.n22 GND 0.153713f
C149 Vout.n23 GND 0.155413f
C150 Vout.t4 GND 0.032704f
C151 Vout.t21 GND 0.032704f
C152 Vout.n24 GND 0.153713f
C153 Vout.n25 GND 0.156222f
C154 Vout.t8 GND 0.032704f
C155 Vout.t20 GND 0.032704f
C156 Vout.n26 GND 0.153713f
C157 Vout.n27 GND 0.210399f
C158 Vout.n28 GND 0.127845f
C159 Vout.n29 GND 0.302213f
C160 Vin.t11 GND 0.33124f
C161 Vin.t14 GND 0.325425f
C162 Vin.n0 GND 0.822091f
C163 Vin.t3 GND 0.041646f
C164 Vin.t9 GND 0.041646f
C165 Vin.n1 GND 0.22387f
C166 Vin.n2 GND 0.523903f
C167 Vin.t17 GND 0.041646f
C168 Vin.t18 GND 0.041646f
C169 Vin.n3 GND 0.228065f
C170 Vin.n4 GND 0.498593f
C171 Vin.t13 GND 0.041646f
C172 Vin.t0 GND 0.041646f
C173 Vin.n5 GND 0.227874f
C174 Vin.n6 GND 0.494534f
C175 Vin.t12 GND 0.041646f
C176 Vin.t4 GND 0.041646f
C177 Vin.n7 GND 0.22515f
C178 Vin.n8 GND 0.395003f
C179 Vin.t6 GND 0.33153f
C180 Vin.t1 GND 0.321965f
C181 Vin.n9 GND 1.00157f
C182 Vin.t2 GND 0.041646f
C183 Vin.t16 GND 0.041646f
C184 Vin.n10 GND 0.229216f
C185 Vin.n11 GND 0.532355f
C186 Vin.t7 GND 0.041646f
C187 Vin.t10 GND 0.041646f
C188 Vin.n12 GND 0.223712f
C189 Vin.n13 GND 0.484973f
C190 Vin.t19 GND 0.041646f
C191 Vin.t15 GND 0.041646f
C192 Vin.n14 GND 0.228449f
C193 Vin.n15 GND 0.491923f
C194 Vin.t5 GND 0.041646f
C195 Vin.t8 GND 0.041646f
C196 Vin.n16 GND 0.22515f
C197 Vin.n17 GND 0.147647f
C198 a_n2515_0.n0 GND 0.946236f
C199 a_n2515_0.t1 GND 0.259367f
C200 a_n2515_0.t3 GND 0.245043f
C201 a_n2515_0.t8 GND 0.245043f
C202 a_n2515_0.t7 GND 0.245043f
C203 a_n2515_0.t0 GND 0.245046f
C204 a_n2515_0.t5 GND 0.242739f
C205 a_n2515_0.t4 GND 0.242739f
C206 a_n2515_0.t2 GND 0.242739f
C207 a_n2515_0.t6 GND 0.242739f
C208 a_n2515_0.t9 GND 0.261642f
C209 a_n2515_0.n1 GND 1.64496f
C210 a_n2515_0.n2 GND 2.08094f
C211 a_n2515_0.n3 GND 0.499303f
C212 a_n2515_0.n4 GND 1.53607f
C213 a_n2515_0.t28 GND 0.061123f
C214 a_n2515_0.t20 GND 0.061123f
C215 a_n2515_0.t12 GND 0.061123f
C216 a_n2515_0.t29 GND 0.060988f
C217 a_n2515_0.t14 GND 0.06089f
C218 a_n2515_0.t21 GND 0.06089f
C219 a_n2515_0.t13 GND 0.06089f
C220 a_n2515_0.t16 GND 0.06089f
C221 a_n2515_0.t22 GND 0.06089f
C222 a_n2515_0.t23 GND 0.06089f
C223 a_n2515_0.t17 GND 0.06089f
C224 a_n2515_0.t25 GND 0.06089f
C225 a_n2515_0.t27 GND 0.06089f
C226 a_n2515_0.t15 GND 0.061123f
C227 a_n2515_0.t26 GND 0.061123f
C228 a_n2515_0.t10 GND 0.061123f
C229 a_n2515_0.t19 GND 0.061123f
C230 a_n2515_0.t18 GND 0.061244f
C231 a_n2515_0.t24 GND 0.061123f
C232 a_n2515_0.t11 GND 0.061123f
.ends

