* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt TOP VINP VOUTP VOUTN VINN CLK VDD VSS
X0 a_478_1100 CLK.t0 VDD.t4 VDD.t3 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X1 VSS CLK.t1 a_304_0 VSS.t3 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X2 VSS a_478_1100 a_2054_0 VSS.t11 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X3 VSS VOUTN.t3 VOUTP.t1 VSS.t6 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X4 VDD a_1207_1100 a_3981_0 VDD.t10 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X5 VDD CLK.t2 a_1207_1100 VDD.t0 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X6 a_3981_0 VOUTP.t3 VOUTN.t1 VDD.t9 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X7 VSS VOUTP.t4 VOUTN.t0 VSS.t0 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X8 a_2054_0 VOUTN.t4 VOUTP.t0 VDD.t8 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X9 VDD a_478_1100 a_2054_0 VDD.t5 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X10 a_478_1100 VINP.t0 a_304_0 VSS.t14 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X11 VOUTP a_478_1100 VSS.t10 VSS.t9 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X12 VOUTN a_1207_1100 VSS.t19 VSS.t18 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X13 a_304_0 VINN.t0 a_1207_1100 VSS.t15 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X14 VSS a_1207_1100 a_3981_0 VSS.t16 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
R0 CLK.n0 CLK.t1 57.2435
R1 CLK CLK.t2 56.5427
R2 CLK.n0 CLK.t0 56.3817
R3 CLK CLK.n0 0.0111579
R4 VDD.n0 VDD.t9 316.795
R5 VDD.n0 VDD.t10 316.195
R6 VDD.n3 VDD.t8 316.195
R7 VDD.n4 VDD.t5 316.195
R8 VDD.n10 VDD.t3 311.132
R9 VDD.n8 VDD.t0 311.132
R10 VDD.n2 VDD.n1 7.15247
R11 VDD.n6 VDD.n5 7.15247
R12 VDD.n9 VDD.n8 2.38511
R13 VDD.n11 VDD.n10 2.38294
R14 VDD.n10 VDD.t4 2.0905
R15 VDD.n8 VDD.n7 2.0905
R16 VDD.n11 VDD.n9 1.33294
R17 VDD.n3 VDD.n2 1.27204
R18 VDD.n9 VDD.n6 0.91974
R19 VDD.n4 VDD.n3 0.6005
R20 VDD.n2 VDD.n0 0.0755
R21 VDD.n6 VDD.n4 0.0755
R22 VDD VDD.n11 0.0449939
R23 VSS.n19 VSS.n18 35712.1
R24 VSS.n45 VSS.n2 32211.3
R25 VSS.n20 VSS.n19 23286.4
R26 VSS.n20 VSS.n2 23286.4
R27 VSS.n23 VSS.n19 13163.2
R28 VSS.n21 VSS.n20 12425.6
R29 VSS.n40 VSS.n2 12267
R30 VSS.n18 VSS.t0 1443.29
R31 VSS.t6 VSS.n21 1443.29
R32 VSS.t14 VSS.t3 989.019
R33 VSS.n41 VSS.n40 812.5
R34 VSS.n40 VSS.t11 726.837
R35 VSS.n44 VSS.t15 716.455
R36 VSS.t16 VSS.n23 706.071
R37 VSS VSS.t14 656.345
R38 VSS.t0 VSS.n17 651.043
R39 VSS.t18 VSS.n10 648.962
R40 VSS.n24 VSS.t16 648.962
R41 VSS.n22 VSS.t6 648.962
R42 VSS.t9 VSS.n4 648.962
R43 VSS.t11 VSS.n39 648.962
R44 VSS.n41 VSS.t15 648.962
R45 VSS.n24 VSS.n10 482.827
R46 VSS.n39 VSS.n4 482.827
R47 VSS.n45 VSS.n44 462.062
R48 VSS.n23 VSS.n22 407.548
R49 VSS.t3 VSS.n45 186.901
R50 VSS.n18 VSS.t18 15.5756
R51 VSS.n21 VSS.t9 15.5756
R52 VSS.n1 VSS.n0 7.11997
R53 VSS.n44 VSS.n43 7.03997
R54 VSS.n42 VSS.n41 7.03997
R55 VSS.n37 VSS.n3 4.50077
R56 VSS.n28 VSS.n27 4.50077
R57 VSS.n32 VSS.n31 4.50063
R58 VSS.n15 VSS.n14 4.50063
R59 VSS.n12 VSS.n11 4.5005
R60 VSS.n9 VSS.n8 4.5005
R61 VSS.n33 VSS.n5 4.5005
R62 VSS.n35 VSS.n34 4.5005
R63 VSS.n17 VSS.n15 3.32886
R64 VSS.n29 VSS.n7 2.3648
R65 VSS.n17 VSS.n16 2.1605
R66 VSS.n37 VSS.n36 2.1605
R67 VSS.n31 VSS.t10 2.1605
R68 VSS.n7 VSS.n6 2.1605
R69 VSS.n27 VSS.n26 2.1605
R70 VSS.n14 VSS.t19 2.1605
R71 VSS.n13 VSS.n10 2.0805
R72 VSS.n25 VSS.n24 2.0805
R73 VSS.n22 VSS.n7 2.0805
R74 VSS.n30 VSS.n4 2.0805
R75 VSS.n39 VSS.n38 2.0805
R76 VSS.n32 VSS.n29 0.965567
R77 VSS.n42 VSS.n3 0.79569
R78 VSS.n29 VSS.n28 0.686453
R79 VSS.n43 VSS.n42 0.59974
R80 VSS VSS.n1 0.485247
R81 VSS.n11 VSS.n8 0.203285
R82 VSS.n34 VSS.n33 0.203285
R83 VSS.n15 VSS.n11 0.166829
R84 VSS.n28 VSS.n8 0.166829
R85 VSS.n33 VSS.n32 0.166829
R86 VSS.n34 VSS.n3 0.166829
R87 VSS.n43 VSS.n1 0.157715
R88 VSS.n35 VSS.n5 0.0244732
R89 VSS.n12 VSS.n9 0.0244732
R90 VSS.n31 VSS.n30 0.0195179
R91 VSS.n38 VSS.n37 0.0195179
R92 VSS.n14 VSS.n13 0.0195179
R93 VSS.n27 VSS.n25 0.0195179
R94 VSS.n30 VSS.n5 0.00103571
R95 VSS.n13 VSS.n12 0.00103571
R96 VSS.n38 VSS.n35 0.000901786
R97 VSS.n25 VSS.n9 0.000901786
R98 VOUTN.n2 VOUTN.t4 56.1724
R99 VOUTN.n2 VOUTN.t3 56.1724
R100 VOUTN.n3 VOUTN.n2 29.048
R101 VOUTN VOUTN.t1 2.56188
R102 VOUTN.n1 VOUTN.n0 2.22447
R103 VOUTN.n1 VOUTN.t0 2.16087
R104 VOUTN.n3 VOUTN.n1 0.3671
R105 VOUTN VOUTN.n3 0.1823
R106 VOUTP VOUTP.t3 56.18
R107 VOUTP.n3 VOUTP.t4 56.0684
R108 VOUTP.n3 VOUTP.n2 20.2978
R109 VOUTP.n2 VOUTP.t0 2.85168
R110 VOUTP.n1 VOUTP.n0 2.22447
R111 VOUTP.n1 VOUTP.t1 2.16087
R112 VOUTP.n2 VOUTP.n1 0.2591
R113 VOUTP VOUTP.n3 0.0969286
R114 VINP VINP.t0 55.9767
R115 VINN VINN.t0 55.9826
C0 CLK VINP 0.014669f
C1 VOUTP VOUTN 1.94745f
C2 a_478_1100 VINP 0.166342f
C3 CLK VINN 0.012448f
C4 a_3981_0 a_1207_1100 0.300768f
C5 VDD a_2054_0 1.24134f
C6 CLK a_1207_1100 0.199918f
C7 VOUTN a_2054_0 0.061728f
C8 VDD a_304_0 0.020392f
C9 VOUTP a_1207_1100 0.201462f
C10 a_478_1100 a_1207_1100 0.232376f
C11 VOUTP a_3981_0 0.163525f
C12 VINP a_304_0 0.037052f
C13 VOUTN VDD 0.589365f
C14 a_304_0 VINN 0.034714f
C15 a_478_1100 CLK 0.324384f
C16 a_478_1100 VOUTP 0.054541f
C17 a_1207_1100 a_2054_0 0.396654f
C18 a_3981_0 a_2054_0 0.089356f
C19 a_1207_1100 a_304_0 0.194884f
C20 a_1207_1100 VDD 0.647286f
C21 a_3981_0 VDD 1.16619f
C22 a_1207_1100 VOUTN 0.198878f
C23 a_3981_0 VOUTN 0.473173f
C24 VOUTP a_2054_0 0.312702f
C25 CLK a_304_0 0.038179f
C26 a_478_1100 a_2054_0 0.229771f
C27 CLK VDD 0.869452f
C28 a_478_1100 a_304_0 0.465024f
C29 a_1207_1100 VINN 0.180516f
C30 VOUTP VDD 0.589635f
C31 a_478_1100 VDD 0.519463f
C32 VINN VSS 0.210259f
C33 VINP VSS 0.2139f
C34 VOUTP VSS 1.69512f
C35 VOUTN VSS 1.66369f
C36 CLK VSS 0.800486f
C37 VDD VSS 12.6574f
C38 a_304_0 VSS 2.25744f
C39 a_3981_0 VSS 0.965151f
C40 a_2054_0 VSS 0.746958f
C41 a_1207_1100 VSS 1.91674f
C42 a_478_1100 VSS 1.71161f
.ends

