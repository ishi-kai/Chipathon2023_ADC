** sch_path: /media/tomoakitanaka/Documents/MyDocuments/personal/ISHIKAI/2024/Chipathon2023_ADC/gitefu/TOP/TOP.sch
.subckt TOP VDD CLK VINP VINN VSS VOUTP VOUTN
*.PININFO VDD:I CLK:I VINP:I VINN:I VSS:I VOUTP:O VOUTN:O
XM1 net3 CLK VSS VSS nfet_03v3 L=0.28u W=2.80u nf=1 m=1
XM2 net1 VINP net3 VSS nfet_03v3 L=0.28u W=2.80u nf=1 m=1
XM4 net1 CLK VDD VDD pfet_03v3 L=0.28u W=2.80u nf=1 m=1
XM6 net4 net1 VDD VDD pfet_03v3 L=0.28u W=2.80u nf=1 m=1
XM7 VOUTP VOUTN net4 VDD pfet_03v3 L=0.28u W=2.80u nf=1 m=1
XM8 net4 net1 VSS VSS nfet_03v3 L=0.28u W=2.80u nf=1 m=1
XM9 VOUTP net1 VSS VSS nfet_03v3 L=0.28u W=2.80u nf=1 m=1
XM10 VOUTP VOUTN VSS VSS nfet_03v3 L=0.28u W=2.80u nf=1 m=1
XM3 net2 VINN net3 VSS nfet_03v3 L=0.28u W=2.80u nf=1 m=1
XM5 net2 CLK VDD VDD pfet_03v3 L=0.28u W=2.80u nf=1 m=1
XM11 net5 net2 VDD VDD pfet_03v3 L=0.28u W=2.80u nf=1 m=1
XM12 VOUTN VOUTP net5 VDD pfet_03v3 L=0.28u W=2.80u nf=1 m=1
XM13 net5 net2 VSS VSS nfet_03v3 L=0.28u W=2.80u nf=1 m=1
XM14 VOUTN net2 VSS VSS nfet_03v3 L=0.28u W=2.80u nf=1 m=1
XM15 VOUTN VOUTP VSS VSS nfet_03v3 L=0.28u W=2.80u nf=1 m=1
.ends
.end
