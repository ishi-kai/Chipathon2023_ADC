* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt TOP VDD CLK VOUTP VOUTN VINP VINN VSS
X0 a_546_n560 VINN.t0 a_n1608_n2000 VSS.t7 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X1 a_546_n560 CLK.t0 VDD.t10 VDD.t9 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X2 VSS a_n1272_n560 a_1616_n2000 VSS.t13 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X3 a_n1608_n2000 CLK.t1 VSS.t6 VSS.t5 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X4 VOUTN a_546_n560 VSS.t4 VSS.t3 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X5 VDD a_n1272_n560 a_1616_n2000 VDD.t3 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X6 VSS a_n1272_n560 VOUTP.t0 VSS.t10 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X7 VOUTP VOUTN.t3 a_1616_n2000 VDD.t2 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X8 a_5710_n560 VOUTP.t3 VOUTN.t2 VDD.t11 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X9 VDD CLK.t2 a_n1272_n560 VDD.t6 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X10 VSS VOUTP.t4 VOUTN.t1 VSS.t16 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X11 a_n1608_n2000 VINP.t0 a_n1272_n560 VSS.t0 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X12 VOUTP VOUTN.t4 VSS.t9 VSS.t8 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X13 a_5710_n560 a_546_n560 VSS.t2 VSS.t1 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X14 a_5710_n560 a_546_n560 VDD.t1 VDD.t0 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
R0 VINN VINN.t0 55.9885
R1 VSS.n24 VSS.n23 11412.8
R2 VSS.n10 VSS.n8 8358.95
R3 VSS.n20 VSS.n19 5254.46
R4 VSS.n24 VSS.n22 5113.97
R5 VSS.n25 VSS.n21 4917.06
R6 VSS.n25 VSS.n24 4917.06
R7 VSS.n9 VSS.n8 4817.7
R8 VSS.n28 VSS.n21 4185.17
R9 VSS.n20 VSS.n8 3516.86
R10 VSS.n21 VSS.n20 3516.86
R11 VSS.n22 VSS.n2 1607.81
R12 VSS.n29 VSS.n28 1510.43
R13 VSS.t3 VSS.n12 1489.42
R14 VSS.t10 VSS.n26 1489.42
R15 VSS.t0 VSS.n0 1489.42
R16 VSS.n18 VSS.n9 1296.56
R17 VSS.n25 VSS.t7 1287.02
R18 VSS.n19 VSS.t16 1088.43
R19 VSS.n19 VSS.t8 989.13
R20 VSS.t13 VSS.n25 569.037
R21 VSS.n13 VSS.n9 551.851
R22 VSS.n28 VSS.n27 517.48
R23 VSS.n13 VSS.t3 477.38
R24 VSS.t16 VSS.n18 477.38
R25 VSS.n29 VSS.t8 477.38
R26 VSS.n27 VSS.t10 477.38
R27 VSS.n26 VSS.t13 477.38
R28 VSS.t7 VSS.n2 477.38
R29 VSS.n1 VSS.t0 477.38
R30 VSS.n23 VSS.n0 418.185
R31 VSS.n12 VSS.n10 402.909
R32 VSS.n22 VSS.n1 110.752
R33 VSS.n10 VSS.t1 74.4717
R34 VSS.n23 VSS.t5 59.1956
R35 VSS.n34 VSS.n2 7.4193
R36 VSS.n36 VSS.n0 7.344
R37 VSS.n35 VSS.n1 7.25447
R38 VSS.n11 VSS.n5 6.1295
R39 VSS VSS.n36 5.1755
R40 VSS.n33 VSS.n4 5.0621
R41 VSS.n32 VSS.n31 4.8875
R42 VSS.n15 VSS.n5 4.8875
R43 VSS.n32 VSS.n5 2.8805
R44 VSS VSS.t6 2.64366
R45 VSS.n7 VSS.n6 2.50972
R46 VSS.n30 VSS.t9 2.50972
R47 VSS.n17 VSS.n16 2.50972
R48 VSS.n14 VSS.t4 2.50972
R49 VSS.n4 VSS.n3 2.45409
R50 VSS.n11 VSS.t2 2.38597
R51 VSS.n12 VSS.n11 2.36672
R52 VSS.n27 VSS.n7 2.26997
R53 VSS.n30 VSS.n29 2.26997
R54 VSS.n18 VSS.n17 2.26997
R55 VSS.n14 VSS.n13 2.26997
R56 VSS.n26 VSS.n4 2.24629
R57 VSS.n34 VSS.n33 1.7285
R58 VSS.n36 VSS.n35 0.9185
R59 VSS.n31 VSS.n30 0.9095
R60 VSS.n33 VSS.n32 0.9005
R61 VSS.n17 VSS.n15 0.7925
R62 VSS.n35 VSS.n34 0.4145
R63 VSS.n15 VSS.n14 0.185
R64 VSS.n31 VSS.n7 0.17375
R65 CLK.n0 CLK.t0 56.8971
R66 CLK.n0 CLK.t2 56.5155
R67 CLK CLK.t1 56.1555
R68 CLK CLK.n0 10.2191
R69 VDD.n7 VDD.t11 322.95
R70 VDD.n8 VDD.t2 321.339
R71 VDD.n5 VDD.t0 311.322
R72 VDD.n4 VDD.t3 311.322
R73 VDD.n0 VDD.t9 311.204
R74 VDD.n2 VDD.t6 311.204
R75 VDD.n9 VDD.n8 11.4455
R76 VDD.n7 VDD.n6 9.7025
R77 VDD.n5 VDD.t1 2.44422
R78 VDD.n4 VDD.n3 2.44422
R79 VDD.n0 VDD.t10 2.23455
R80 VDD.n2 VDD.n1 2.23455
R81 VDD.n8 VDD.n7 2.1905
R82 VDD.n6 VDD.n5 0.635
R83 VDD.n6 VDD.n4 0.4865
R84 VDD.n9 VDD.n2 0.2535
R85 VDD VDD.n0 0.1705
R86 VDD VDD.n9 0.1355
R87 VOUTN.n3 VOUTN.t3 68.0895
R88 VOUTN VOUTN.t4 56.0655
R89 VOUTN.n3 VOUTN.n2 9.7565
R90 VOUTN VOUTN.n3 9.2165
R91 VOUTN.n1 VOUTN.n0 3.55417
R92 VOUTN.n1 VOUTN.t2 3.32705
R93 VOUTN.n2 VOUTN.t1 3.09022
R94 VOUTN.n2 VOUTN.n1 1.2245
R95 VOUTP.n4 VOUTP.t3 67.9167
R96 VOUTP VOUTP.t4 56.0475
R97 VOUTP.n4 VOUTP.n3 9.7565
R98 VOUTP VOUTP.n4 9.1175
R99 VOUTP.n1 VOUTP.t0 3.69547
R100 VOUTP.n1 VOUTP.n0 3.12815
R101 VOUTP.n3 VOUTP.n2 2.88322
R102 VOUTP.n3 VOUTP.n1 1.535
R103 VINP VINP.t0 55.9885
C0 VINP a_n1272_n560 0.077845f
C1 CLK a_n1272_n560 0.454491f
C2 a_1616_n2000 a_n1272_n560 0.278387f
C3 VOUTP VOUTN 1.22218f
C4 VOUTN a_546_n560 0.828295f
C5 VOUTP a_546_n560 0.380564f
C6 CLK VDD 0.793055f
C7 a_5710_n560 VDD 1.02449f
C8 VINN a_546_n560 0.042096f
C9 VDD a_n1272_n560 0.530103f
C10 VDD a_1616_n2000 1.03301f
C11 a_n1608_n2000 a_546_n560 0.175682f
C12 VINN a_n1608_n2000 0.025074f
C13 a_5710_n560 VOUTN 0.256955f
C14 VOUTN a_n1272_n560 0.305764f
C15 a_5710_n560 VOUTP 0.133657f
C16 a_1616_n2000 VOUTN 0.141823f
C17 VOUTP a_n1272_n560 0.695778f
C18 CLK a_546_n560 0.045468f
C19 a_5710_n560 a_546_n560 0.728923f
C20 a_n1272_n560 a_546_n560 0.193251f
C21 a_1616_n2000 VOUTP 0.277948f
C22 a_1616_n2000 a_546_n560 0.64116f
C23 VINN a_n1272_n560 0.012743f
C24 a_n1608_n2000 VINP 0.037779f
C25 VDD VOUTN 0.576678f
C26 VDD VOUTP 0.615516f
C27 CLK a_n1608_n2000 0.044894f
C28 VDD a_546_n560 1.73142f
C29 a_n1608_n2000 a_n1272_n560 0.274203f
C30 VINN VSS 0.229258f
C31 VINP VSS 0.218379f
C32 VOUTP VSS 3.43853f
C33 VOUTN VSS 3.55699f
C34 CLK VSS 1.36602f
C35 VDD VSS 15.025001f
C36 a_n1608_n2000 VSS 3.24777f
C37 a_5710_n560 VSS 2.14206f
C38 a_1616_n2000 VSS 1.99211f
C39 a_546_n560 VSS 5.04437f
C40 a_n1272_n560 VSS 3.00793f
.ends

