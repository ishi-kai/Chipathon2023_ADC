* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt TOP VDD CLK VOUTP VOUTN VINP VINN VSS
X0 a_546_n560 VINN.t0 a_n1608_n2000 VSS.t9 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X1 a_546_n560 CLK.t0 VDD.t10 VDD.t9 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X2 VSS a_n1272_n560 a_1616_n2000 VSS.t14 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X3 a_n1608_n2000 CLK.t1 VSS.t8 VSS.t7 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X4 VOUTN a_546_n560 VSS.t6 VSS.t5 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X5 VDD a_n1272_n560 a_1616_n2000 VDD.t3 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X6 VSS a_n1272_n560 VOUTP.t2 VSS.t11 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X7 VOUTP VOUTN.t3 a_1616_n2000 VDD.t11 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X8 a_5710_n560 VOUTP.t3 VOUTN.t2 VDD.t2 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X9 VDD CLK.t2 a_n1272_n560 VDD.t6 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X10 VSS VOUTP.t4 VOUTN.t0 VSS.t0 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X11 a_n1608_n2000 VINP.t0 a_n1272_n560 VSS.t10 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X12 VOUTP VOUTN.t4 VSS.t18 VSS.t17 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X13 a_5710_n560 a_546_n560 VSS.t4 VSS.t3 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X14 a_5710_n560 a_546_n560 VDD.t1 VDD.t0 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
R0 VINN VINN.t0 55.9885
R1 VSS.n24 VSS.n23 11412.8
R2 VSS.n10 VSS.n8 8358.95
R3 VSS.n20 VSS.n19 5254.46
R4 VSS.n24 VSS.n22 5113.97
R5 VSS.n25 VSS.n21 4917.06
R6 VSS.n25 VSS.n24 4917.06
R7 VSS.n9 VSS.n8 4817.7
R8 VSS.n28 VSS.n21 4185.17
R9 VSS.n20 VSS.n8 3516.86
R10 VSS.n21 VSS.n20 3516.86
R11 VSS.n22 VSS.n2 1607.81
R12 VSS.n29 VSS.n28 1510.43
R13 VSS.t5 VSS.n12 1489.42
R14 VSS.t11 VSS.n26 1489.42
R15 VSS.t10 VSS.n0 1489.42
R16 VSS.n18 VSS.n9 1296.56
R17 VSS.n25 VSS.t9 1287.02
R18 VSS.n19 VSS.t0 1088.43
R19 VSS.n19 VSS.t17 989.13
R20 VSS.t14 VSS.n25 569.037
R21 VSS.n13 VSS.n9 551.851
R22 VSS.n28 VSS.n27 517.48
R23 VSS.n13 VSS.t5 477.38
R24 VSS.t0 VSS.n18 477.38
R25 VSS.n29 VSS.t17 477.38
R26 VSS.n27 VSS.t11 477.38
R27 VSS.n26 VSS.t14 477.38
R28 VSS.t9 VSS.n2 477.38
R29 VSS.n1 VSS.t10 477.38
R30 VSS.n23 VSS.n0 418.185
R31 VSS.n12 VSS.n10 402.909
R32 VSS.n22 VSS.n1 110.752
R33 VSS.n10 VSS.t3 74.4717
R34 VSS.n23 VSS.t7 59.1956
R35 VSS.n34 VSS.n2 7.4193
R36 VSS.n36 VSS.n0 7.344
R37 VSS.n35 VSS.n1 7.25447
R38 VSS.n11 VSS.n5 6.1295
R39 VSS VSS.n36 5.1755
R40 VSS.n33 VSS.n4 5.0621
R41 VSS.n32 VSS.n31 4.8875
R42 VSS.n15 VSS.n5 4.8875
R43 VSS.n32 VSS.n5 2.8805
R44 VSS VSS.t8 2.64366
R45 VSS.n7 VSS.n6 2.50972
R46 VSS.n30 VSS.t18 2.50972
R47 VSS.n17 VSS.n16 2.50972
R48 VSS.n14 VSS.t6 2.50972
R49 VSS.n4 VSS.n3 2.45409
R50 VSS.n11 VSS.t4 2.38597
R51 VSS.n12 VSS.n11 2.36672
R52 VSS.n27 VSS.n7 2.26997
R53 VSS.n30 VSS.n29 2.26997
R54 VSS.n18 VSS.n17 2.26997
R55 VSS.n14 VSS.n13 2.26997
R56 VSS.n26 VSS.n4 2.24629
R57 VSS.n34 VSS.n33 1.7285
R58 VSS.n36 VSS.n35 0.9185
R59 VSS.n31 VSS.n30 0.9095
R60 VSS.n33 VSS.n32 0.9005
R61 VSS.n17 VSS.n15 0.7925
R62 VSS.n35 VSS.n34 0.4145
R63 VSS.n15 VSS.n14 0.185
R64 VSS.n31 VSS.n7 0.17375
R65 CLK.n0 CLK.t0 56.8971
R66 CLK.n0 CLK.t2 56.5155
R67 CLK CLK.t1 56.1555
R68 CLK CLK.n0 10.2191
R69 VDD.n7 VDD.t2 322.95
R70 VDD.n8 VDD.t11 321.339
R71 VDD.n5 VDD.t0 311.322
R72 VDD.n4 VDD.t3 311.322
R73 VDD.n0 VDD.t9 311.204
R74 VDD.n2 VDD.t6 311.204
R75 VDD.n9 VDD.n8 11.4455
R76 VDD.n7 VDD.n6 9.7025
R77 VDD.n5 VDD.t1 2.44422
R78 VDD.n4 VDD.n3 2.44422
R79 VDD.n0 VDD.t10 2.23455
R80 VDD.n2 VDD.n1 2.23455
R81 VDD.n8 VDD.n7 2.1905
R82 VDD.n6 VDD.n5 0.635
R83 VDD.n6 VDD.n4 0.4865
R84 VDD.n9 VDD.n2 0.2535
R85 VDD VDD.n0 0.1705
R86 VDD VDD.n9 0.1355
R87 VOUTN.n3 VOUTN.t3 68.0895
R88 VOUTN VOUTN.t4 56.0655
R89 VOUTN.n3 VOUTN.n2 9.7565
R90 VOUTN VOUTN.n3 9.2165
R91 VOUTN.n1 VOUTN.n0 3.55417
R92 VOUTN.n1 VOUTN.t2 3.32705
R93 VOUTN.n2 VOUTN.t0 3.09022
R94 VOUTN.n2 VOUTN.n1 1.2245
R95 VOUTP.n4 VOUTP.t3 67.9167
R96 VOUTP VOUTP.t4 56.0475
R97 VOUTP.n4 VOUTP.n3 9.7565
R98 VOUTP VOUTP.n4 9.1175
R99 VOUTP.n1 VOUTP.t2 3.69547
R100 VOUTP.n1 VOUTP.n0 3.12815
R101 VOUTP.n3 VOUTP.n2 2.88322
R102 VOUTP.n3 VOUTP.n1 1.535
R103 VINP VINP.t0 55.9885
C0 VOUTN w_2022_n798 0.017717f
C1 a_1616_n2000 a_n1272_n560 0.278387f
C2 a_5710_n560 a_546_n560 0.728923f
C3 VDD a_546_n560 1.73142f
C4 VOUTP w_6672_n798 0.017717f
C5 w_n24_n798 CLK 0.017949f
C6 a_546_n560 a_n1608_n2000 0.175682f
C7 VOUTN a_n1272_n560 0.305764f
C8 VOUTP a_546_n560 0.380564f
C9 VDD a_5710_n560 1.02449f
C10 VINP a_n1272_n560 0.077845f
C11 VOUTN a_1616_n2000 0.141823f
C12 VOUTP a_5710_n560 0.133657f
C13 VINN a_546_n560 0.042096f
C14 VOUTP VDD 0.615516f
C15 a_546_n560 CLK 0.045468f
C16 VINN a_n1608_n2000 0.025074f
C17 VDD CLK 0.793055f
C18 CLK a_n1608_n2000 0.044894f
C19 a_n1272_n560 w_3674_n798 0.017717f
C20 w_5140_n800 a_546_n560 0.017877f
C21 a_n1272_n560 a_546_n560 0.193251f
C22 a_1616_n2000 a_546_n560 0.64116f
C23 a_n1272_n560 VDD 0.530103f
C24 w_n1510_n798 CLK 0.017949f
C25 a_n1272_n560 a_n1608_n2000 0.274203f
C26 a_1616_n2000 VDD 1.03301f
C27 a_n1272_n560 VOUTP 0.695778f
C28 VOUTN a_546_n560 0.828295f
C29 VOUTN a_5710_n560 0.256955f
C30 a_n1272_n560 VINN 0.012743f
C31 a_1616_n2000 VOUTP 0.277948f
C32 VOUTN VDD 0.576678f
C33 a_n1272_n560 CLK 0.454491f
C34 VOUTN VOUTP 1.22218f
C35 VINP a_n1608_n2000 0.037779f
C36 VINN VSS 0.228664f
C37 VINP VSS 0.217057f
C38 VOUTP VSS 3.42015f
C39 VOUTN VSS 3.53867f
C40 CLK VSS 1.33f
C41 VDD VSS 15.025001f
C42 a_n1608_n2000 VSS 3.24777f
C43 a_5710_n560 VSS 2.14206f
C44 a_1616_n2000 VSS 1.99211f
C45 a_546_n560 VSS 5.0256f
C46 a_n1272_n560 VSS 2.98937f
.ends

