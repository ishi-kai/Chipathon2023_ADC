* NGSPICE file created from SAR_TOP.ext - technology: gf180mcuD

.subckt SAR_TOP VIN VSS VDD XRST CLK OUT[1] OUT[0] OUT[3] OUT[2] OUT[5] OUT[4] EOC
X0 VDD.t1021 a_41180_n2804 a_41092_n2760 VDD.t1020 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1 a_23932_n20052 a_23844_n20008 VSS.t1943 VSS.t1942 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2 a_32533_n14520 a_32413_n14564 a_31789_n14564 VSS.t1657 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X3 a_46556_n2804 a_46468_n2760 VSS.t1266 VSS.t1265 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4 VDD.t1333 a_47452_n16916 a_47364_n16872 VDD.t1332 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X5 a_11087_n7460.t29 a_11023_n6840.t20 a_13501_n6460.t11 VDD.t107 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X6 a_46108_n12212 a_46020_n12168 VSS.t4244 VSS.t4243 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7 VSS.t1647 a_24233_n13388 a_24128_n13248 VSS.t1646 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X8 VSS.t984 a_28764_n8247 a_30228_n8203 VSS.t983 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X9 VDD.t3641 a_47452_n13780 a_47364_n13736 VDD.t3640 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X10 VDD.t1296 a_30396_n7508 a_30240_n7464 VDD.t1295 pfet_06v0 ad=0.4392p pd=1.94u as=0.4758p ps=2u w=1.22u l=0.5u
X11 VSS.t429 a_21772_n8292.t8 a_13623_n17552.t7 VSS.t428 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X12 a_46780_n20485 a_46692_n20388 VSS.t4230 VSS.t4229 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X13 VSS.t55 a_11023_n14874.t20 a_11087_n15494.t29 VSS.t54 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X14 VDD.t3525 a_40060_n7508 a_39972_n7464 VDD.t3524 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X15 VDD.t411 a_28721_n9076.t2 a_30324_n10600 VDD.t410 pfet_06v0 ad=0.4005p pd=2.12u as=0.1456p ps=1.08u w=0.56u l=0.5u
X16 VDD.t2056 a_33564_n20052 a_33476_n20008 VDD.t1162 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X17 VDD.t4226 a_45212_n16916 a_45124_n16872 VDD.t4225 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X18 a_38716_n9076 a_38628_n9032 VSS.t1617 VSS.t1616 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X19 VDD.t4228 a_45212_n13780 a_45124_n13736 VDD.t4227 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X20 VDD.t1547 a_40060_n4372 a_39972_n4328 VDD.t1546 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X21 a_21692_n5468.t7 a_26440_n5940.t4 VSS.t399 VSS.t398 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X22 VDD.t936 a_43084_n18917 a_42996_n18820 VDD.t935 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X23 a_11087_n18172.t29 a_11023_n17552.t20 VSS.t410 VSS.t58 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X24 a_38403_n5503 a_38733_n5431 a_38853_n5874 VDD.t2165 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X25 VSS.t1333 a_32560_n7020 a_32455_n7420 VSS.t1332 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
D0 VSS.t191 a_26388_n17606.t2 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X26 VDD.t1864 a_31324_n20052 a_31236_n20008 VDD.t1863 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X27 a_44540_n20485 a_44452_n20388 VSS.t4250 VSS.t4249 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X28 a_43420_n20485 a_43332_n20388 VSS.t1624 VSS.t1623 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X29 a_32668_n16916 a_32580_n16872 VSS.t2138 VSS.t2137 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X30 VSS.t373 a_10778_2852.t15 a_10712_4516.t19 VSS.t372 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X31 VSS.t236 a_44640_1944.t8 OUT[5].t7 VSS.t235 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X32 a_38403_n2367 a_38733_n2295 a_38853_n2738 VDD.t2750 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X33 a_13501_n9138.t19 a_13623_n9518.t8 a_11087_n10138.t26 VSS.t239 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X34 a_47452_n20052 a_47364_n20008 VSS.t978 VSS.t977 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X35 VDD.t1150 a_38716_n18484 a_38628_n18440 VDD.t1149 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X36 a_47004_n5940 a_46916_n5896 VSS.t1444 VSS.t1443 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X37 a_11023_n22908.t9 a_13623_n22908.t8 VSS.t203 VSS.t202 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X38 a_30428_n16916 a_30340_n16872 VSS.t991 VSS.t990 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X39 VDD.t4192 a_37844_1564 a_38256_1564.t7 VDD.t4191 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X40 a_38295_332 a_39056_820 a_38847_464 VSS.t1011 nfet_06v0 ad=0.2007p pd=1.475u as=94.5f ps=0.885u w=0.36u l=0.6u
X41 a_39648_n2020 a_26553_377.t2 VDD.t138 VDD.t137 pfet_06v0 ad=0.2486p pd=2.01u as=0.35315p ps=1.96u w=0.565u l=0.5u
X42 a_31628_n5940.t31 a_33496_n6659.t8 VDD.t158 VDD.t157 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X43 a_45212_n20052 a_45124_n20008 VSS.t2455 VSS.t2454 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X44 VDD.t2154 a_31772_n18484 a_31684_n18440 VDD.t2153 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X45 VDD.t2536 a_34860_n3189 a_34756_n3140 VDD.t2535 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X46 a_25237_n4327 a_24233_n3980 VSS.t1939 VSS.t1938 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X47 a_44428_n9509 a_44340_n9412 VSS.t3618 VSS.t3617 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X48 a_23564_n17700 a_28568_n16066 VSS.t4270 VSS.t4269 nfet_06v0 ad=0.1261p pd=1.005u as=0.2134p ps=1.85u w=0.485u l=0.6u
X49 a_27984_376 a_27884_332.t2 VDD.t692 VDD.t691 pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X50 a_28156_n6412.t7 a_29800_n5940.t7 VSS.t752 VSS.t751 nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X51 VSS.t116 a_11023_n12196.t20 a_11087_n12816.t9 VSS.t54 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X52 VDD.t630 a_21772_n20836.t8 a_13623_n6840.t15 VDD.t629 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X53 a_13623_n6840.t14 a_21772_n20836.t9 VDD.t666 VDD.t665 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X54 a_28645_n13252 a_21692_n6694.t2 a_28437_n13705 VSS.t673 nfet_06v0 ad=0.1722p pd=1.24u as=0.3608p ps=2.52u w=0.82u l=0.6u
X55 a_23212_n12124 a_22904_n12080 VDD.t2242 VDD.t2241 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X56 a_33780_n5112 a_24815_n3588.t4 a_33604_n5112 VSS.t16 nfet_06v0 ad=0.1312p pd=1.14u as=0.1148p ps=1.1u w=0.82u l=0.6u
X57 VDD.t1858 a_43980_n7941 a_43892_n7844 VDD.t1857 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X58 a_30696_n704 a_29856_n1121 a_30408_n1104 VSS.t1007 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X59 VDD.t958 a_43980_n4805 a_43892_n4708 VDD.t957 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X60 a_26736_n364 a_21692_n5468.t16 VSS.t393 VSS.t392 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X61 VSS.t29 a_45648_1564.t8 EOC.t7 VSS.t28 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X62 VDD.t1300 a_42188_n6373 a_42100_n6276 VDD.t1299 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X63 VSS.t3282 a_24681_n7116 a_24576_n6976 VSS.t3281 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X64 a_32262_n452 a_22444_332.t7 VSS.t324 VSS.t323 nfet_06v0 ad=0.3608p pd=2.52u as=0.2911p ps=1.53u w=0.82u l=0.6u
X65 a_32424_n10512 a_31460_n10116 a_32220_n10512 VSS.t1325 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X66 a_11087_n23528.t30 a_2167_3472.t72 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X67 VDD.t2891 a_42188_n3237 a_42100_n3140 VDD.t2890 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X68 a_42748_n9076 a_42660_n9032 VSS.t1327 VSS.t1326 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X69 a_21772_n12996 a_25831_n12996 VDD.t2545 VDD.t2544 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X70 a_33048_n7420 a_32560_n7020 a_33308_n7376 VDD.t1286 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X71 VDD.t2576 a_35356_n16916 a_35268_n16872 VDD.t2575 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X72 a_13623_n4162.t15 a_21772_1116.t4 VDD.t620 VDD.t619 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X73 VDD.t1852 a_22588_n20052 a_22500_n20008 VDD.t1851 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X74 a_36588_n15348 a_36500_n15304 VSS.t4282 VSS.t4212 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X75 VDD.t23 a_24815_n3588.t5 a_23004_n2332 VDD.t22 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X76 a_13501_n9138.t0 a_11023_n9518.t20 a_11087_n10138.t0 VDD.t541 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
D1 VSS.t477 a_23072_n13432.t8 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X77 VSS.t326 a_22444_332.t8 a_33252_n1192 VSS.t325 nfet_06v0 ad=0.2911p pd=1.53u as=0.3608p ps=2.52u w=0.82u l=0.6u
X78 VSS.t646 a_29920_n3900.t2 a_24815_n3588.t0 VSS.t645 nfet_06v0 ad=0.2112p pd=1.84u as=0.1248p ps=1u w=0.48u l=0.6u
X79 VDD.t932 a_33116_n16916 a_33028_n16872 VDD.t931 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X80 a_27605_n8456 a_27485_n8500 a_26861_n8567 VSS.t1016 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X81 a_33564_n20485 a_33476_n20388 VSS.t2136 VSS.t2135 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X82 a_34348_n15348 a_34260_n15304 VSS.t2257 VSS.t2256 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X83 VDD.t572 a_21772_n3588.t4 a_13623_n20230.t15 VDD.t571 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X84 a_34552_n3140 a_34000_n3140 a_34348_n3140 VDD.t2706 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X85 a_21772_n8292.t7 a_23564_n8292 VDD.t1178 VDD.t1177 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X86 a_34232_n2272 a_32432_n2689 a_33292_n2716 VSS.t3471 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X87 VDD.t3523 a_40508_n9076 a_40420_n9032 VDD.t3522 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X88 a_32444_n20485 a_32356_n20388 VSS.t2621 VSS.t2620 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X89 VDD.t4176 a_31451_n7508 a_25020_n8200.t1 VDD.t4175 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X90 a_47564_n4805 a_47476_n4708 VSS.t1611 VSS.t1610 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X91 a_35356_n20052 a_35268_n20008 VSS.t1506 VSS.t1505 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X92 VDD.t1448 a_35244_n15348 a_35156_n15304 VDD.t953 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X93 VSS.t887 a_4001_4292.t3 a_10778_2852.t10 VSS.t342 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X94 a_30204_n20485 a_30116_n20388 VSS.t1382 VSS.t1381 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X95 a_11087_n15494.t19 a_11023_n14874.t21 a_13501_n14494.t19 VDD.t73 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X96 a_34708_n5896.t7 a_33776_n5896.t7 VSS.t872 VSS.t871 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X97 a_30324_n10600 a_29076_n8292.t4 a_30136_n10600 VDD.t439 pfet_06v0 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.5u
X98 VDD.t2435 a_24220_n15260 a_24116_n15216 VDD.t2434 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X99 a_21996_332.t1 a_27884_332.t3 VDD.t694 VDD.t693 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X100 a_33116_n20052 a_33028_n20008 VSS.t4278 VSS.t4277 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X101 a_39500_n3237 a_39412_n3140 VSS.t2238 VSS.t2237 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X102 a_27190_n5112 a_26358_n4618 a_27022_n5112 VSS.t1454 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X103 VSS.t479 a_23072_n13432.t9 a_23024_n10112 VSS.t478 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X104 VDD.t2720 a_33004_n15348 a_32916_n15304 VDD.t2719 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X105 VSS.t1631 a_31965_n8292 a_32085_n8248 VSS.t1630 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X106 a_46220_n12645 a_46132_n12548 VSS.t1615 VSS.t1614 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X107 a_13501_n17172.t19 a_11023_n17552.t21 a_11087_n18172.t19 VDD.t400 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X108 a_10712_4516.t0 a_3935_4156.t3 VSS.t452 VSS.t378 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X109 OUT[1].t15 a_33216_1944.t8 VDD.t421 VDD.t420 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X110 VSS.t431 a_21772_n8292.t9 a_13623_n17552.t6 VSS.t430 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X111 a_26172_n18484 a_26084_n18440 VSS.t997 VSS.t996 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X112 a_11087_n18172.t18 a_11023_n17552.t22 a_13501_n17172.t18 VDD.t401 pfet_03v3 ad=0.728p pd=3.32u as=1.82p ps=6.9u w=2.8u l=0.28u
X113 VDD.t1397 a_34895_n1192 a_35351_n1170 VDD.t1396 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X114 a_21772_n11428.t7 a_23564_n11428 VDD.t1671 VDD.t1670 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X115 a_25472_n14816 a_23360_n15233 a_25160_n14816 VDD.t1454 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X116 a_34403_332 a_34068_n4 VDD.t1856 VDD.t1855 pfet_06v0 ad=0.3477p pd=1.79u as=0.4392p ps=1.94u w=1.22u l=0.5u
X117 a_32100_n1976 a_29076_n8292.t5 a_32308_n1976 VSS.t466 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X118 VDD.t1553 a_35800_n3456 a_36217_n3500 VDD.t1552 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X119 a_32856_n7376 a_32455_n7420 a_31799_n7508 VSS.t4320 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X120 VDD.t1790 a_47564_n11077 a_47476_n10980 VDD.t1789 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X121 a_39724_n17349 a_39636_n17252 VSS.t1984 VSS.t1983 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X122 a_27301_n16388 a_21692_n6694.t3 VSS.t675 VSS.t674 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X123 a_31548_n10172.t7 a_33496_n8222.t7 VSS.t292 VSS.t291 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X124 a_39724_n14213 a_39636_n14116 VSS.t3715 VSS.t3714 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X125 OUT[5].t6 a_44640_1944.t9 VSS.t238 VSS.t237 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X126 VDD.t4162 a_47900_n1236 a_47812_n1192 VDD.t2657 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X127 VDD.t970 a_40620_n5940 a_40532_n5896 VDD.t969 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X128 VDD.t978 a_45324_n11077 a_45236_n10980 VDD.t977 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X129 VSS.t2130 a_26635_n12996 a_26547_n12951 VSS.t2129 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X130 a_47452_n5940 a_47364_n5896 VSS.t1260 VSS.t1259 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X131 a_11087_n12816.t19 a_11023_n12196.t21 a_13501_n11816.t9 VDD.t127 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X132 VDD.t928 a_43196_n18484 a_43108_n18440 VDD.t927 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X133 a_31660_n17349 a_31572_n17252 VSS.t2953 VSS.t2952 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X134 VDD.t3649 a_33467_1116 a_30732_332.t1 VDD.t3648 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X135 a_25020_n11383 a_28721_n9076.t3 VSS.t421 VSS.t420 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X136 VDD.t1587 a_21772_n452.t4 a_13623_n22908.t0 VDD.t1586 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X137 VDD.t2441 a_47004_n1669 a_46916_n1572 VDD.t2440 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X138 VSS.t4226 a_34652_n11391 a_34350_n10980 VSS.t4225 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X139 a_25612_n878.t1 a_27259_804.t2 a_36709_n2276 VSS.t849 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X140 VDD.t2354 a_31656_n704 a_32073_n844 VDD.t2353 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X141 a_26915_n2672 a_25895_n2624 VDD.t3633 VDD.t3632 pfet_06v0 ad=0.101p pd=0.905u as=0.3975p ps=2.185u w=0.505u l=0.5u
X142 a_27093_n8248 a_26973_n8292 VSS.t1026 VSS.t1025 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X143 a_44876_n9509 a_44788_n9412 VSS.t2445 VSS.t2444 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X144 a_28009_n12168 a_27279_n12146 VDD.t2551 VDD.t2550 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X145 a_28868_n9387 a_28519_n10160.t2 a_28624_n9394 VDD.t786 pfet_06v0 ad=0.58035p pd=2.155u as=0.4012p ps=1.85u w=1.095u l=0.5u
X146 a_25237_n13735 a_24233_n13388 VDD.t1572 VDD.t1571 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X147 VDD.t160 a_33496_n6659.t9 a_31628_n5940.t30 VDD.t159 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X148 VSS.t3005 a_26643_n8292 a_23887_n5156 VSS.t3004 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X149 a_28437_n13705 a_22220_690.t2 VDD.t776 VDD.t775 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X150 VSS.t888 a_4001_4292.t4 a_10778_2852.t11 VSS.t344 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X151 OUT[3].t15 a_38256_1564.t8 VDD.t190 VDD.t189 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X152 VDD.t4157 a_46220_n17349 a_46132_n17252 VDD.t4156 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X153 a_23524_464 a_23404_816 VDD.t1564 VDD.t1563 pfet_06v0 ad=0.1313p pd=1.025u as=0.22725p ps=1.91u w=0.505u l=0.5u
X154 a_43532_n3237 a_43444_n3140 VSS.t1195 VSS.t1194 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X155 VDD.t2234 a_24684_n16432 a_22600_n12124 VDD.t2233 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X156 a_13623_n20230.t7 a_21772_n3588.t5 VSS.t608 VSS.t607 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X157 a_23360_n11680 a_23212_n12124 a_23192_n11680 VSS.t2617 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X158 VDD.t4172 a_46220_n14213 a_46132_n14116 VDD.t4171 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X159 a_24693_n6680 a_24573_n6724 a_23949_n6724 VSS.t2630 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X160 a_36364_n12645 a_36276_n12548 VSS.t1457 VSS.t1456 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X161 VSS.t45 a_21692_n5111.t2 a_24628_n363 VSS.t44 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X162 a_30988_n18917 a_30900_n18820 VSS.t1233 VSS.t1232 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X163 a_11087_n23528.t13 a_11023_n22908.t20 a_13501_n22528.t19 VDD.t206 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X164 a_42771_769 a_43101_841 a_43221_951 VSS.t1929 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X165 a_34124_n12645 a_34036_n12548 VSS.t2006 VSS.t2005 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X166 a_29868_n17349 a_29780_n17252 VSS.t1178 VSS.t1177 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D2 VSS.t327 a_22444_332.t9 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X167 VSS.t375 a_10778_2852.t16 a_10712_4516.t18 VSS.t374 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X168 VDD.t1133 a_36588_n11077 a_36500_n10980 VDD.t1132 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X169 VSS.t764 a_24481_761.t8 a_26115_n328 VSS.t763 nfet_06v0 ad=0.1224p pd=1.04u as=0.134p ps=1.1u w=0.36u l=0.6u
X170 VDD.t1271 a_44509_n452 a_44629_168 VDD.t1270 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X171 a_21692_n13308.t7 a_26328_n6654.t7 VSS.t2661 VSS.t2660 nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X172 a_28736_n4633.t13 a_30452_n5156.t3 VDD.t1039 VDD.t1038 pfet_06v0 ad=0.2197p pd=1.365u as=0.4056p ps=1.805u w=0.845u l=0.5u
X173 VSS.t1502 a_26531_n8639 a_22712_n7420 VSS.t1501 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X174 VDD.t1131 a_40956_n9076 a_40868_n9032 VDD.t1130 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X175 a_40956_n13780 a_40868_n13736 VSS.t968 VSS.t967 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X176 a_26123_n1976 a_25647_n1976 VSS.t1998 VSS.t1997 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X177 VDD.t3516 a_43084_n9509 a_42996_n9412 VDD.t3515 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X178 VDD.t1129 a_25084_1564 a_33216_1944.t7 VDD.t1128 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X179 a_46108_n7508 a_46020_n7464 VSS.t1498 VSS.t1497 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X180 a_40956_n10644 a_40868_n10600 VSS.t1424 VSS.t1423 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D3 a_22220_690.t3 VDD.t777 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X181 VDD.t3118 a_46220_n7941 a_46132_n7844 VDD.t3117 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X182 a_31856_n11296 a_29332_n11301 a_31544_n11296 VSS.t3560 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X183 a_38716_n12212 a_38628_n12168 VSS.t3236 VSS.t3235 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X184 VDD.t3376 a_27736_1248 a_28153_1204 VDD.t3375 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X185 VDD.t3571 a_27167_n10808 a_27623_n10830 VDD.t3570 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X186 VDD.t2889 a_46220_n4805 a_46132_n4708 VDD.t2888 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X187 VSS.t4157 a_35456_n4628.t7 a_32108_n2332.t7 VSS.t4156 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X188 a_23479_n5156 a_26943_n7442 VSS.t2951 VSS.t2950 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X189 VDD.t4108 a_25940_n17606.t2 a_21772_n9860 VDD.t4107 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X190 VDD.t3428 a_37820_n16916 a_37732_n16872 VDD.t3427 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X191 a_25831_n12996 a_27526_n13714 VDD.t2232 VDD.t2231 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X192 a_32499_n3844 a_32359_n4372 a_31787_n3969 VSS.t2596 nfet_06v0 ad=0.217p pd=1.515u as=0.3586p ps=2.51u w=0.815u l=0.6u
X193 VSS.t1305 a_24752_n8292 a_22140_n6694.t0 VSS.t1304 nfet_06v0 ad=0.2344p pd=1.56u as=0.3608p ps=2.52u w=0.82u l=0.6u
X194 a_30820_n3544 a_29920_n3900.t3 a_30616_n3544 VSS.t647 nfet_06v0 ad=0.1722p pd=1.24u as=0.1722p ps=1.24u w=0.82u l=0.6u
X195 a_33497_n9032 a_32767_n9010 VDD.t1119 VDD.t1118 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X196 a_21692_n18917 a_21604_n18820 VSS.t1165 VSS.t1164 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X197 VDD.t4104 a_36700_n16916 a_36612_n16872 VDD.t4103 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X198 VDD.t1738 a_37820_n13780 a_37732_n13736 VDD.t1737 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X199 VDD.t905 a_35692_n18917 a_35604_n18820 VDD.t904 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X200 VDD.t2423 a_37484_n17349 a_37396_n17252 VDD.t2422 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X201 a_30040_n3844 a_29920_n3900.t4 a_29846_n3844 VSS.t648 nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X202 a_26551_n7464 a_26095_n7464 VDD.t1115 VDD.t1114 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X203 VDD.t1206 a_23932_n20052 a_23844_n20008 VDD.t1205 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X204 a_31544_1248 a_29744_1564 a_30604_1515 VSS.t1158 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X205 VDD.t2521 a_37484_n14213 a_37396_n14116 VDD.t2520 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X206 a_32100_n1976 a_32860_n2020 VSS.t3604 VSS.t3603 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X207 a_22672_n2214.t0 a_21916_n1975 VSS.t1156 VSS.t1155 nfet_06v0 ad=0.2569p pd=1.56u as=0.2244p ps=1.9u w=0.51u l=0.6u
X208 a_30599_n12167 a_30871_n11728 a_30787_n12167 VDD.t897 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X209 VDD.t702 a_24481_761.t9 a_33868_n4240 VDD.t701 pfet_06v0 ad=0.45p pd=2.02u as=0.3432p ps=2.44u w=0.78u l=0.5u
X210 VDD.t2517 a_33452_n18917 a_33364_n18820 VDD.t2516 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X211 VDD.t1434 a_35244_n17349 a_35156_n17252 VDD.t1433 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D4 a_24481_761.t10 VDD.t703 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X212 VDD.t1106 a_32332_n18917 a_32244_n18820 VDD.t1105 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X213 a_43084_n17349 a_42996_n17252 VSS.t955 VSS.t954 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X214 VDD.t1369 a_35244_n14213 a_35156_n14116 VDD.t1368 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X215 a_30296_1564 a_29332_1243 a_30092_1564 VSS.t2589 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X216 a_32449_n704 a_23072_n13432.t10 VSS.t481 VSS.t480 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X217 a_30584_n1954 a_29444_n4328.t6 VDD.t1496 VDD.t1495 pfet_06v0 ad=0.4488p pd=2.92u as=0.458p ps=2.02u w=1.02u l=0.5u
X218 VDD.t1831 a_23619_n6724 a_22264_n5852 VDD.t1830 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X219 a_24609_n13248 a_23072_n13432.t11 VSS.t483 VSS.t482 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X220 VDD.t1524 a_38268_n7508 a_38180_n7464 VDD.t1523 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X221 a_37820_n20052 a_37732_n20008 VSS.t1294 VSS.t1293 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X222 a_43084_n14213 a_42996_n14116 VSS.t3650 VSS.t3649 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X223 VDD.t3029 a_29900_760.t2 a_29812_860 VDD.t3028 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X224 VDD.t1514 a_27988_n4328 a_31348_n1931 VDD.t1513 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X225 VSS.t568 a_13623_n4162.t16 a_11023_n4162.t9 VSS.t567 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X226 VDD.t1511 a_46556_n10644 a_46468_n10600 VDD.t1510 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X227 a_36700_n20052 a_36612_n20008 VSS.t1290 VSS.t1289 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X228 a_42476_1515 a_42168_1564 VDD.t1721 VDD.t1720 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X229 VDD.t1503 a_47452_n1669 a_47364_n1572 VDD.t1502 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X230 a_26630_n5112 a_26154_n4536 a_26358_n4618 VSS.t1961 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X231 a_23108_n12080 a_23072_n13432.t12 VDD.t462 VDD.t461 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X232 a_26098_n9240 a_25642_n9816 VDD.t2235 VDD.t996 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X233 VDD.t1560 a_47452_n20052 a_47364_n20008 VDD.t1559 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X234 a_11087_n20850.t30 a_2167_3472.t15 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X235 a_30555_n13780 a_30903_n13780 VDD.t2504 VDD.t2503 pfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X236 a_27175_860 a_24815_n3588.t6 a_26991_860 VSS.t17 nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X237 a_27829_n15512 a_27709_n16132 a_27085_n16132 VDD.t3503 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X238 VDD.t632 a_21692_n6694.t4 a_28437_n13705 VDD.t631 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X239 a_37785_n364 a_24481_761.t11 VDD.t705 VDD.t704 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X240 a_25936_1564 a_25524_1243 VDD.t1367 VDD.t1366 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X241 VDD.t2230 a_48012_n101 a_47924_n4 VDD.t2023 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X242 a_41653_n1170 a_41533_n727 VDD.t3548 VDD.t3547 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X243 a_22220_n9860 a_24492_n5156 a_24388_n4708 VDD.t3498 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X244 VDD.t1148 a_45212_n20052 a_45124_n20008 VDD.t1147 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X245 a_47452_1900 a_47364_1944 VSS.t938 VSS.t937 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X246 VSS.t1414 a_28492_332 a_28444_860 VSS.t1413 nfet_06v0 ad=0.2132p pd=1.34u as=98.399994f ps=1.06u w=0.82u l=0.6u
X247 VDD.t2229 a_39612_n4805 a_39524_n4708 VDD.t2228 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X248 a_46556_n16916 a_46468_n16872 VSS.t3628 VSS.t3627 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X249 VDD.t140 a_31628_n5940.t32 a_29800_n5940.t6 VDD.t139 pfet_06v0 ad=0.3608p pd=2.52u as=0.2952p ps=1.54u w=0.82u l=0.5u
X250 VDD.t879 a_32413_n12996 a_32533_n12376 VDD.t878 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X251 VDD.t1357 a_27804_n14165 a_27700_n14116 VDD.t1356 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X252 a_11023_n6840.t0 a_13623_n6840.t16 VSS.t718 VSS.t717 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X253 a_46668_n6373 a_46580_n6276 VSS.t1135 VSS.t1134 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X254 a_24368_n14816 a_24220_n15260 a_24200_n14816 VSS.t2519 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X255 a_43980_n3237 a_43892_n3140 VSS.t3952 VSS.t3951 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X256 VDD.t3372 a_45660_n18484 a_45572_n18440 VDD.t3371 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X257 VDD.t2281 a_30192_n15304.t7 a_24481_761.t0 VDD.t1642 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X258 VDD.t4019 a_42476_1515 a_42372_1564 VDD.t4018 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X259 a_27055_n1192 a_26431_n1192 a_26907_n616 VSS.t3278 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X260 a_11087_n12816.t30 a_2167_3472.t30 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X261 VSS.t1043 a_21772_n17700.t8 a_13623_n9518.t0 VSS.t1042 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X262 a_23072_n13432.t0 a_29744_n15604.t7 VDD.t1637 VDD.t1636 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X263 a_11087_n7460.t28 a_11023_n6840.t21 a_13501_n6460.t10 VDD.t108 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X264 VDD.t3868 a_44540_n18484 a_44452_n18440 VDD.t3867 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X265 a_13623_n9518.t1 a_21772_n17700.t9 VSS.t1045 VSS.t1044 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X266 VSS.t1851 a_21772_n14564.t4 a_13623_n12196.t7 VSS.t1850 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X267 a_22672_n2214.t1 a_22820_n2804 a_22672_n2759 VDD.t3866 pfet_06v0 ad=0.3159p pd=1.735u as=0.44955p ps=1.955u w=1.215u l=0.5u
X268 a_22856_n10112 a_22016_n10529 a_22568_n10512 VSS.t1955 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X269 VSS.t927 a_40652_n1572 a_45648_1564.t3 VSS.t926 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X270 a_27032_51 a_26736_n364 a_25975_n184 VDD.t1470 pfet_06v0 ad=0.2424p pd=1.465u as=0.25375p ps=1.51u w=0.505u l=0.5u
X271 a_33496_n6659.t0 CLK.t0 VSS.t1013 VSS.t1012 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X272 a_28841_n8548 a_28721_n9076.t4 a_28617_n8548 VSS.t422 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X273 a_13623_n12196.t6 a_21772_n14564.t5 VSS.t2080 VSS.t2079 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X274 VDD.t4058 a_22140_n6694.t2 a_27281_n16854 VDD.t4057 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X275 VDD.t1414 a_31760_n12168 a_33280_n13248 VDD.t1413 pfet_06v0 ad=0.3432p pd=2.44u as=0.2028p ps=1.3u w=0.78u l=0.5u
X276 VDD.t1872 a_33832_n8572 a_25612_n6679 VDD.t1871 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X277 a_28624_n9394 a_24348_n16087.t2 VDD.t2425 VDD.t2424 pfet_06v0 ad=0.4012p pd=1.85u as=0.4972p ps=3.14u w=1.13u l=0.5u
X278 VDD.t1344 a_42300_n18484 a_42212_n18440 VDD.t1343 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X279 VSS.t1949 a_22164_n2760 a_28841_n3844 VSS.t1948 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X280 a_29920_n3900.t0 a_31787_n3969 VSS.t1597 VSS.t1596 nfet_06v0 ad=0.2119p pd=1.335u as=0.3586p ps=2.51u w=0.815u l=0.6u
X281 a_29560_n3544 a_29920_n3900.t5 a_31248_n3544 VSS.t649 nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X282 a_47116_n9509 a_47028_n9412 VSS.t1397 VSS.t1396 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X283 a_21692_n13308.t6 a_26328_n6654.t8 VSS.t2663 VSS.t2662 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X284 a_27964_n20052 a_27876_n20008 VSS.t1030 VSS.t1029 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X285 a_35324_1564 a_34872_1619 VDD.t1408 VDD.t1407 pfet_06v0 ad=0.2028p pd=1.3u as=0.45p ps=2.02u w=0.78u l=0.5u
X286 VSS.t557 a_11023_n9518.t21 a_11087_n10138.t1 VSS.t68 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X287 VSS.t190 a_26388_n17606.t3 a_22220_690.t0 VSS.t189 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X288 VSS.t1345 a_13623_n14874.t16 a_11023_n14874.t0 VSS.t1344 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X289 EOC.t15 a_45648_1564.t9 VDD.t46 VDD.t45 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X290 OUT[2].t15 a_37024_1944.t8 VDD.t1687 VDD.t1686 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X291 VSS.t1448 a_32262_n452 a_25940_n17606.t0 VSS.t1447 nfet_06v0 ad=0.2911p pd=1.53u as=0.2132p ps=1.34u w=0.82u l=0.6u
X292 a_21692_n13308.t15 a_26328_n6654.t9 VDD.t2607 VDD.t2606 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X293 a_46556_n7508 a_46468_n7464 VSS.t1395 VSS.t1394 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X294 a_30787_n12167 a_30871_n11728 a_30807_n11684 VSS.t959 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X295 a_25724_n20052 a_25636_n20008 VSS.t1393 VSS.t1392 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X296 a_11023_n14874.t1 a_13623_n14874.t17 VSS.t1347 VSS.t1346 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X297 a_26047_n4328 a_25423_n4328 a_25879_n4328 VDD.t1336 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X298 a_43196_n12212 a_43108_n12168 VSS.t1663 VSS.t1662 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X299 VSS.t1922 a_11023_n20230.t20 a_11087_n20850.t0 VSS.t60 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X300 VSS.t4159 a_35456_n4628.t8 a_32108_n2332.t6 VSS.t4158 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X301 a_27302_n13160 a_26470_n13736 a_27154_n13736 VDD.t1211 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X302 a_24573_n12996 a_21872_n12530 VDD.t1868 VDD.t1867 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X303 VSS.t75 a_13623_n17552.t16 a_11023_n17552.t9 VSS.t74 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X304 a_42076_n2804 a_41988_n2760 VSS.t1386 VSS.t1385 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X305 VDD.t1462 a_35356_n20052 a_35268_n20008 VDD.t1461 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X306 VDD.t3964 a_47004_n16916 a_46916_n16872 VDD.t3963 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X307 a_26643_n8292 a_26973_n8292 a_27093_n8248 VSS.t1024 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X308 VDD.t3924 a_47004_n13780 a_46916_n13736 VDD.t3923 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X309 a_25860_n9032 a_25412_n8501 VSS.t1484 VSS.t1483 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X310 a_28433_n8548 a_25573_n12167 VSS.t2174 VSS.t2173 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X311 VDD.t2049 a_33116_n20052 a_33028_n20008 VDD.t2048 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X312 a_46332_n20485 a_46244_n20388 VSS.t3593 VSS.t3592 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X313 VDD.t1422 a_40060_n16916 a_39972_n16872 VDD.t1421 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X314 OUT[1].t14 a_33216_1944.t9 VDD.t423 VDD.t422 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X315 a_11087_n7460.t19 a_11023_n6840.t22 VSS.t104 VSS.t56 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X316 VDD.t1719 a_37932_n11077 a_37844_n10980 VDD.t1718 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X317 VSS.t1814 a_31664_n13292 a_31559_n13692 VSS.t1813 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X318 a_32736_n1572 a_32636_n2020 a_32308_n1976 VDD.t876 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X319 VDD.t3977 a_40060_n13780 a_39972_n13736 VDD.t3976 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X320 a_1955_4292.t1 a_2167_3472.t84 a_n199_2852 VSS.t330 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X321 VDD.t598 a_29920_n3900.t6 a_29444_n4328.t3 VDD.t597 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X322 VDD.t688 a_29800_n5940.t8 a_28156_n6412.t15 VDD.t687 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X323 VSS.t1581 a_34089_n10252 a_33984_n10112 VSS.t1580 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X324 VSS.t1821 a_13623_n12196.t16 a_11023_n12196.t0 VSS.t1820 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X325 VDD.t2333 a_24236_2258.t2 a_22444_2253.t7 VDD.t2332 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X326 a_37680_n320 a_35568_n4 a_37368_n320 VDD.t4014 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
D5 a_10712_4516.t30 VDD.t324 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X327 VSS.t766 a_24481_761.t12 a_38435_864 VSS.t765 nfet_06v0 ad=0.1224p pd=1.04u as=0.134p ps=1.1u w=0.36u l=0.6u
X328 VDD.t707 a_24481_761.t13 a_31787_n3969 VDD.t706 pfet_06v0 ad=0.33755p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X329 a_11023_n12196.t1 a_13623_n12196.t17 VSS.t1823 VSS.t1822 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X330 a_31011_n8292 a_31341_n8292 a_31461_n7694 VDD.t3975 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X331 a_47004_n20052 a_46916_n20008 VSS.t1699 VSS.t1698 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X332 VDD.t1104 a_33564_n18484 a_33476_n18440 VDD.t1103 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X333 VDD.t2609 a_26328_n6654.t10 a_21692_n13308.t14 VDD.t2608 pfet_06v0 ad=0.367p pd=1.92u as=0.4392p ps=1.94u w=1.22u l=0.5u
X334 VSS.t677 a_21692_n6694.t5 a_30532_n8548 VSS.t676 nfet_06v0 ad=0.3608p pd=2.52u as=0.1148p ps=1.1u w=0.82u l=0.6u
X335 a_32158_n12212 a_31961_n11340 VDD.t4010 VDD.t4009 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X336 a_27960_n320 a_27032_51 a_27792_n320 VSS.t919 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X337 VDD.t1615 a_26383_n2968 a_26839_n2990 VDD.t1614 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X338 VSS.t1571 a_27744_n12908 a_27639_n12537 VSS.t1570 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X339 VDD.t2091 a_31324_n18484 a_31236_n18440 VDD.t2090 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X340 a_26383_1944 a_25759_1944 a_26215_1944 VDD.t892 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X341 a_40060_n20052 a_39972_n20008 VSS.t1708 VSS.t1707 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X342 a_21772_n20836.t7 a_23564_n20836 VDD.t889 VDD.t888 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X343 a_27700_n14116 a_26532_n14437 a_27496_n14116 VDD.t1962 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X344 a_33272_n2272 a_32432_n2689 a_32984_n2672 VSS.t3470 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X345 a_24945_n11680 a_23072_n13432.t13 VSS.t485 VSS.t484 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X346 a_27224_n62 a_26631_7 a_27960_n320 VSS.t1488 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
D6 a_21692_n6694.t6 VDD.t633 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X347 a_10778_2852.t11 a_4001_4292.t5 VSS.t889 VSS.t346 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X348 a_11023_n20230.t9 a_13623_n20230.t16 VSS.t614 VSS.t613 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X349 a_42277_n1192 a_42157_n660 a_41533_n727 VDD.t1711 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X350 a_35064_n11383 a_34350_n10980 VSS.t1520 VSS.t1519 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X351 VSS.t616 a_13623_n20230.t17 a_11023_n20230.t8 VSS.t615 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X352 VDD.t1725 a_38268_n16916 a_38180_n16872 VDD.t1724 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X353 a_33280_n13248 a_31559_n13692 a_32152_n13692 VDD.t3991 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X354 a_24233_n3980 a_23072_n13432.t14 VDD.t464 VDD.t463 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X355 a_28624_n9394 a_27281_n16854 a_28644_n9815 VSS.t1989 nfet_06v0 ad=0.3586p pd=2.51u as=0.2119p ps=1.335u w=0.815u l=0.6u
X356 a_27281_n16854 a_21692_n6694.t7 VDD.t635 VDD.t634 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X357 VSS.t3979 a_29408_1944.t8 OUT[0].t7 VSS.t3978 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X358 VDD.t2051 a_29532_n4372.t4 a_29444_n4328.t4 VDD.t2050 pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X359 VDD.t1733 a_38268_n13780 a_38180_n13736 VDD.t1732 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X360 a_30500_1564 a_24481_761.t14 VDD.t709 VDD.t708 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X361 a_24573_n9860 a_24965_n9860 VSS.t2062 VSS.t2061 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X362 VDD.t3746 a_47900_n10644 a_47812_n10600 VDD.t3745 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X363 a_11023_n22908.t8 a_13623_n22908.t9 VSS.t205 VSS.t204 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X364 a_33496_n6659.t1 CLK.t1 VSS.t1896 VSS.t1895 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X365 a_10712_4516.t17 a_10778_2852.t17 VSS.t377 VSS.t376 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X366 VDD.t873 a_40652_n1572 a_45648_1564.t7 VDD.t872 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X367 VSS.t2750 a_11023_n4162.t20 VSS.t2750 VSS.t58 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.28u
X368 a_22016_n5825 a_21604_n5412 VSS.t3581 VSS.t3580 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X369 a_29908_n6980 a_25612_n6679 VSS.t1277 VSS.t1276 nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X370 a_41404_n7508 a_41316_n7464 VSS.t3808 VSS.t3807 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X371 VDD.t3854 a_39612_n9076 a_39524_n9032 VDD.t3853 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X372 a_35356_n20485 a_35268_n20388 VSS.t3801 VSS.t3800 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X373 VDD.t3063 a_40196_1944 a_41392_1944.t7 VDD.t1781 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X374 a_29920_n3900.t1 a_31787_n3969 VDD.t1532 VDD.t1531 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X375 VDD.t387 a_26440_n5940.t5 a_21692_n5468.t15 VDD.t386 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X376 VDD.t3855 a_24573_n9860 a_24693_n9240 VDD.t996 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X377 a_38268_n20052 a_38180_n20008 VSS.t3150 VSS.t3149 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X378 a_47564_n9509 a_47476_n9412 VSS.t3938 VSS.t3937 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X379 a_33116_n20485 a_33028_n20388 VSS.t3799 VSS.t3798 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X380 a_24088_n16087 a_24348_n16087.t3 VDD.t2427 VDD.t2426 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X381 a_47900_n16916 a_47812_n16872 VSS.t3551 VSS.t3550 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X382 a_42244_n1572 a_29900_760.t3 a_42096_n1572 VDD.t3030 pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X383 a_44316_n1669 a_44228_n1572 VSS.t3505 VSS.t3504 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X384 a_13501_n19850.t19 a_13623_n20230.t18 a_11087_n20850.t29 VSS.t617 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X385 VDD.t3852 a_22588_n18484 a_22500_n18440 VDD.t1239 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X386 VSS.t3129 a_33533_908 a_33653_952 VSS.t3128 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
D7 a_22444_332.t10 VDD.t317 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X387 a_33984_n10112 a_31460_n10116 a_33672_n10112 VSS.t1324 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X388 a_43084_n4805 a_42996_n4708 VSS.t3930 VSS.t3929 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X389 a_21692_n13308.t13 a_26328_n6654.t11 VDD.t2611 VDD.t2610 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X390 a_44876_n18917 a_44788_n18820 VSS.t3934 VSS.t3933 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X391 VDD.t2283 a_30192_n15304.t8 a_24481_761.t1 VDD.t2282 pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X392 a_30192_n15304.t6 a_27988_n20388 VDD.t2739 VDD.t715 pfet_06v0 ad=0.2952p pd=1.54u as=0.3608p ps=2.52u w=0.82u l=0.5u
X393 a_48012_n12645 a_47924_n12548 VSS.t3503 VSS.t3502 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X394 a_22876_n13692 a_22568_n13648 VSS.t3875 VSS.t3874 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X395 a_46220_n3237 a_46132_n3140 VSS.t3548 VSS.t3547 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X396 a_42636_n18917 a_42548_n18820 VSS.t3873 VSS.t3872 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X397 a_n263_3472.t15 a_22444_2253.t8 VDD.t2336 VDD.t451 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X398 a_26266_n9240 a_25642_n9816 a_26098_n9240 VDD.t996 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X399 VDD.t1055 a_28972_n17349 a_28884_n17252 VDD.t1054 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X400 a_36812_n7941 a_36724_n7844 VSS.t1480 VSS.t1479 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X401 a_21916_n6694.t1 a_33494_n9860 VDD.t1053 VDD.t1052 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X402 a_44092_n4372 a_44004_n4328 VSS.t1565 VSS.t1564 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X403 VDD.t4008 a_31961_n11340 a_31856_n11296 VDD.t4007 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X404 a_35692_n17349 a_35604_n17252 VSS.t3925 VSS.t3924 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X405 a_43644_n705 a_43833_1204 VDD.t3416 VDD.t3415 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X406 VSS.t2840 a_39357_n2228 a_39477_n2184 VSS.t2839 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X407 a_32108_n2332.t5 a_35456_n4628.t9 VSS.t4161 VSS.t4160 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X408 VDD.t3790 a_47900_n5940 a_47812_n5896 VDD.t3789 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X409 a_28132_376 a_22444_332.t11 a_27984_376 VDD.t318 pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X410 a_46693_951 a_46573_841 VSS.t2807 VSS.t2806 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X411 VDD.t2730 a_47116_n11077 a_47028_n10980 VDD.t2729 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X412 a_35692_n14213 a_35604_n14116 VSS.t3537 VSS.t2248 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X413 VDD.t2760 a_47900_n2804 a_47812_n2760 VDD.t2759 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X414 a_33452_n17349 a_33364_n17252 VSS.t2836 VSS.t2835 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X415 VDD.t458 a_21772_1116.t5 a_13623_n4162.t14 VDD.t457 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X416 a_37820_n7508 a_37732_n7464 VSS.t3869 VSS.t3868 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X417 VDD.t3687 a_41292_n11077 a_41204_n10980 VDD.t3686 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X418 a_26215_n2968 a_25759_n3544 VDD.t3483 VDD.t3482 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X419 VDD.t2758 a_40172_n11077 a_40084_n10980 VDD.t2757 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X420 a_30192_n15304.t2 a_27988_n20388 VSS.t2812 VSS.t529 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X421 a_33452_n14213 a_33364_n14116 VSS.t2832 VSS.t2831 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X422 VSS.t768 a_24481_761.t15 a_32499_n3844 VSS.t767 nfet_06v0 ad=0.1224p pd=1.04u as=0.217p ps=1.515u w=0.36u l=0.6u
X423 VSS.t703 a_28156_n6412.t16 a_26328_n6654.t2 VSS.t702 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X424 VDD.t3683 a_43644_n9076 a_43556_n9032 VDD.t3682 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X425 a_45660_n12212 a_45572_n12168 VSS.t3583 VSS.t3582 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X426 a_13501_n22528.t9 a_13623_n22908.t10 a_11087_n23528.t9 VSS.t206 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X427 a_31212_n17349 a_31124_n17252 VSS.t3626 VSS.t3625 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X428 a_35064_1506 a_34471_1575 a_35800_1248 VSS.t4037 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
D8 a_23072_n13432.t15 VDD.t465 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X429 a_44540_n12212 a_44452_n12168 VSS.t4023 VSS.t4022 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D9 VSS.t486 a_23072_n13432.t16 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X430 a_47900_n9076 a_47812_n9032 VSS.t3833 VSS.t3832 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X431 VDD.t3459 a_26266_n9240 a_26702_n9240 VDD.t996 pfet_06v0 ad=0.1656p pd=1.28u as=61.199993f ps=0.7u w=0.36u l=0.5u
X432 VDD.t2243 a_37820_n20052 a_37732_n20008 VDD.t961 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X433 VDD.t2237 a_36700_n20052 a_36612_n20008 VDD.t2236 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X434 a_28144_n4708 a_27414_n5112 VDD.t3845 VDD.t3844 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X435 a_42300_n12212 a_42212_n12168 VSS.t3885 VSS.t3884 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X436 a_32152_n13692 a_31664_n13292 a_32412_n13648 VDD.t1729 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X437 a_21772_n452.t0 a_23564_n452.t2 VDD.t3658 VDD.t3657 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X438 VDD.t3674 a_46220_n18917 a_46132_n18820 VDD.t3673 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X439 VDD.t3450 a_48012_n17349 a_47924_n17252 VDD.t3449 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X440 VSS.t1622 a_34403_332 a_34271_376 VSS.t1621 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X441 VSS.t1718 a_29744_n15604.t8 a_23072_n13432.t1 VSS.t1717 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X442 a_29800_n9815 a_28624_n9394 VDD.t4210 VDD.t4209 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X443 a_35804_n16916 a_35716_n16872 VSS.t3485 VSS.t3484 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X444 VDD.t3050 a_48012_n14213 a_47924_n14116 VDD.t3049 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X445 a_23072_n13432.t2 a_29744_n15604.t9 VSS.t1720 VSS.t1719 nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
D10 a_23072_n13432.t17 VDD.t466 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X446 VSS.t453 a_3935_4156.t4 a_10712_4516.t1 VSS.t380 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X447 a_34708_n5896.t15 a_33776_n5896.t8 VDD.t828 VDD.t827 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X448 VDD.t1815 CLK.t2 a_33496_n6659.t2 VDD.t1814 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X449 a_38156_n12645 a_38068_n12548 VSS.t3146 VSS.t3145 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X450 VDD.t4217 a_23816_n13248 a_24233_n13388 VDD.t4216 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X451 a_22856_n8544 a_22016_n8961 a_22568_n8944 VSS.t3866 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X452 OUT[1].t7 a_33216_1944.t10 VSS.t437 VSS.t436 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X453 a_37632_n2020 a_36388_n1572 VDD.t1032 VDD.t1031 pfet_06v0 ad=0.2486p pd=2.01u as=0.35315p ps=1.96u w=0.565u l=0.5u
D11 VSS.t678 a_21692_n6694.t8 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X454 a_22772_n1104 a_23072_n13432.t18 VDD.t468 VDD.t467 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X455 VSS.t1890 a_37585_n3140 a_38171_n3544 VSS.t1889 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X456 a_22856_n5408 a_22016_n5825 a_22568_n5808 VSS.t3152 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X457 a_23220_n7376 a_22052_n6980 a_23016_n7376 VDD.t1492 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X458 VDD.t3445 a_33999_n1400 a_34455_n1422 VDD.t3444 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X459 a_28736_1944 a_22500_n1976 VSS.t1794 VSS.t1793 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X460 a_24716_n5156.t1 a_24233_n8684 VDD.t1024 VDD.t415 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X461 a_40956_n18484 a_40868_n18440 VSS.t1551 VSS.t1550 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X462 a_21804_n2273.t0 a_32132_2428 VSS.t3483 VSS.t3482 nfet_06v0 ad=0.3608p pd=2.52u as=0.2344p ps=1.56u w=0.82u l=0.6u
X463 VDD.t2756 a_40732_n2804 a_40644_n2760 VDD.t2755 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X464 a_41852_n7508 a_41764_n7464 VSS.t3479 VSS.t3478 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X465 a_13501_n9138.t1 a_11023_n9518.t22 a_11087_n10138.t2 VDD.t542 pfet_03v3 ad=1.82p pd=6.9u as=0.728p ps=3.32u w=2.8u l=0.28u
X466 a_40956_n15348 a_40868_n15304 VSS.t2830 VSS.t2829 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X467 a_42748_n13780 a_42660_n13736 VSS.t1549 VSS.t1548 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X468 a_25237_n13735 a_24233_n13388 VSS.t1645 VSS.t1644 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X469 a_29295_n1400 a_28671_n1976 a_29147_n1976 VSS.t3864 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X470 VDD.t389 a_26440_n5940.t6 a_21692_n5468.t14 VDD.t388 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X471 a_33815_1384 a_34471_1575 a_34367_1619 VDD.t3958 pfet_06v0 ad=0.25375p pd=1.51u as=0.1313p ps=1.025u w=0.505u l=0.5u
X472 a_25237_n10599 a_24233_n10252 VSS.t1038 VSS.t1037 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X473 a_42748_n10644 a_42660_n10600 VSS.t1540 VSS.t1539 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X474 a_30808_n6334 a_30215_n6265 a_31544_n6592 VSS.t1888 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X475 a_44764_n1669 a_44676_n1572 VSS.t1769 VSS.t1768 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X476 VDD.t1678 a_23816_n8544 a_24233_n8684 VDD.t513 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X477 a_40508_n13780 a_40420_n13736 VSS.t1884 VSS.t1883 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X478 a_40508_n10644 a_40420_n10600 VSS.t1886 VSS.t1885 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X479 VDD.t1803 a_41852_n15348 a_41764_n15304 VDD.t1802 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D12 a_24481_761.t16 VDD.t710 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X480 a_24752_n16132 a_24716_n5156.t2 VDD.t1324 VDD.t1323 pfet_06v0 ad=0.2486p pd=2.01u as=0.35315p ps=1.96u w=0.565u l=0.5u
X481 EOC.t14 a_45648_1564.t10 VDD.t48 VDD.t47 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X482 VDD.t1799 a_30740_n7464 a_31936_n6592 VDD.t1798 pfet_06v0 ad=0.3432p pd=2.44u as=0.2028p ps=1.3u w=0.78u l=0.5u
X483 VDD.t1342 a_27964_n20052 a_27876_n20008 VDD.t1341 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X484 VDD.t2486 a_39612_n16916 a_39524_n16872 VDD.t2485 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X485 VDD.t393 a_21692_n5468.t17 a_22724_860.t1 VDD.t392 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X486 a_34392_n9815 a_25972_n6276 VDD.t1797 VDD.t1796 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X487 a_23484_n18917 a_23396_n18820 VSS.t2557 VSS.t2556 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X488 VDD.t1794 a_37484_n18917 a_37396_n18820 VDD.t1793 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X489 VDD.t966 a_39612_n13780 a_39524_n13736 VDD.t965 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D13 VSS.t769 a_24481_761.t17 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X490 VDD.t1217 a_25724_n20052 a_25636_n20008 VDD.t1216 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X491 VDD.t1675 a_39276_n17349 a_39188_n17252 VDD.t1674 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X492 a_37820_n20485 a_37732_n20388 VSS.t1522 VSS.t1521 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X493 VDD.t3529 a_39276_n14213 a_39188_n14116 VDD.t3528 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X494 VDD.t995 a_24233_n10252 a_24128_n10112 VDD.t994 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X495 a_35692_n13780 a_35604_n13736 VSS.t2798 VSS.t2797 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X496 VDD.t3779 a_35244_n18917 a_35156_n18820 VDD.t3778 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X497 VDD.t1786 a_37036_n17349 a_36948_n17252 VDD.t1785 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X498 a_11023_n6840.t1 a_13623_n6840.t17 VSS.t720 VSS.t719 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X499 VDD.t3627 a_37036_n14213 a_36948_n14116 VDD.t3626 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X500 a_39612_n20052 a_39524_n20008 VSS.t1654 VSS.t1653 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X501 a_23212_n12124 a_22904_n12080 VSS.t2317 VSS.t2316 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X502 a_24693_n12952 a_24573_n12996 a_23949_n12996 VSS.t2643 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X503 a_11023_n22908.t19 a_13623_n22908.t11 VDD.t217 VDD.t216 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X504 VDD.t2079 a_32152_n13692 a_31960_n13648 VDD.t2078 pfet_06v0 ad=0.2222p pd=1.89u as=0.2424p ps=1.465u w=0.505u l=0.5u
X505 VDD.t4032 a_23932_n18484 a_23844_n18440 VDD.t3554 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X506 a_34649_n2412 a_24481_761.t18 VDD.t712 VDD.t711 pfet_06v0 ad=0.3159p pd=1.735u as=0.33755p ps=1.955u w=1.215u l=0.5u
X507 VDD.t2041 a_30676_n7844 a_31919_n9032 VDD.t2040 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X508 a_43416_1248 a_41204_1243 a_42476_1515 VDD.t1784 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X509 VSS.t1960 a_26154_n4536 a_26630_n5112 VSS.t1959 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X510 VDD.t2039 a_46108_n10644 a_46020_n10600 VDD.t2038 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X511 a_30604_n11029 a_30296_n10980 VDD.t4031 VDD.t4030 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X512 a_27302_n13160 a_26470_n13736 a_27134_n13160 VSS.t1269 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X513 VSS.t329 a_22444_332.t12 a_27572_860 VSS.t328 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X514 a_31459_n14564 a_31789_n14564 a_31909_n13966 VDD.t2480 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X515 VDD.t917 a_28764_n8247 a_30228_n8203 VDD.t916 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X516 a_24128_n13248 a_21604_n13252 a_23816_n13248 VSS.t2219 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X517 VDD.t1262 a_21804_n2273.t2 a_24516_n14475 VDD.t1261 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X518 VDD.t1516 a_47004_n20052 a_46916_n20008 VDD.t1515 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X519 OUT[1].t13 a_33216_1944.t11 VDD.t425 VDD.t424 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X520 a_34986_n9032 a_29532_n10311 a_34092_n9076 VDD.t3985 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X521 a_34538_n10980 a_22140_n6694.t3 a_34350_n10980 VDD.t4059 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X522 a_24233_n13388 a_23072_n13432.t19 VDD.t470 VDD.t469 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X523 a_21772_1116.t0 a_23564_1116.t2 VDD.t3409 VDD.t2343 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X524 a_40508_n4372 a_40420_n4328 VSS.t2214 VSS.t2213 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X525 VDD.t4017 a_40060_n20052 a_39972_n20008 VDD.t3563 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X526 a_46108_n16916 a_46020_n16872 VSS.t2212 VSS.t2211 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X527 a_23912_n15216 a_22948_n14820 a_23708_n15216 VSS.t2109 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X528 VDD.t2032 a_47004_n7508 a_46916_n7464 VDD.t2031 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X529 a_22164_n2760 a_21716_n2229 VSS.t4080 VSS.t4079 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X530 VDD.t2130 a_47004_n4372 a_46916_n4328 VDD.t2129 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X531 a_25559_n10980 a_25831_n11428 a_24684_n16432 VDD.t1773 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X532 a_11087_n20850.t1 a_11023_n20230.t21 a_13501_n19850.t9 VDD.t1842 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X533 VDD.t4271 a_47452_n18484 a_47364_n18440 VDD.t4270 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X534 a_30903_n13780 a_31559_n13692 a_31455_n13648 VDD.t3990 pfet_06v0 ad=0.25375p pd=1.51u as=0.1313p ps=1.025u w=0.505u l=0.5u
X535 VSS.t651 a_29920_n3900.t7 a_24815_n3588.t1 VSS.t650 nfet_06v0 ad=0.1248p pd=1u as=0.2112p ps=1.84u w=0.48u l=0.6u
X536 a_34708_n5896.t14 a_33776_n5896.t9 VDD.t830 VDD.t829 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X537 a_31628_n5940.t15 a_33496_n6659.t10 VSS.t142 VSS.t141 nfet_06v0 ad=0.1261p pd=1.005u as=0.2134p ps=1.85u w=0.485u l=0.6u
X538 a_42188_n6373 a_42100_n6276 VSS.t1190 VSS.t1189 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X539 a_21772_n17700.t3 a_23564_n17700 VSS.t4312 VSS.t4311 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X540 VDD.t1770 a_28636_n16916 a_28548_n16872 VDD.t1769 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X541 a_34872_1619 a_34576_1204 a_33815_1384 VDD.t1568 pfet_06v0 ad=0.2424p pd=1.465u as=0.25375p ps=1.51u w=0.505u l=0.5u
X542 VDD.t3032 a_29900_760.t4 a_33508_n408 VDD.t3031 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X543 a_42412_n5940 a_42324_n5896 VSS.t2099 VSS.t2098 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X544 VDD.t254 a_13623_n9518.t9 a_11023_n9518.t19 VDD.t253 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X545 VDD.t1187 a_45212_n18484 a_45124_n18440 VDD.t1186 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D14 VSS.t831 a_22220_690.t4 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X546 a_21772_n14564.t0 a_23564_n14564.t2 VSS.t3810 VSS.t3809 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X547 VSS.t241 a_13623_n9518.t10 a_11023_n9518.t9 VSS.t240 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X548 a_26266_n13736 a_25642_n13736 a_26118_n13160 VSS.t1231 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X549 a_48012_332 a_47924_376 VSS.t2097 VSS.t2096 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X550 a_28009_n1192.t0 a_27279_n1170 VSS.t2196 VSS.t2195 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X551 a_34860_n3189 a_34552_n3140 VDD.t1780 VDD.t1779 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X552 a_27628_n18484 a_27540_n18440 VSS.t4335 VSS.t4334 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X553 VDD.t1663 a_21692_n16916 a_21604_n16872 VDD.t1662 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X554 a_32579_769 a_32909_841 a_33029_951 VSS.t4315 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X555 a_11023_n9518.t8 a_13623_n9518.t11 VSS.t243 VSS.t242 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X556 a_21872_n9394 a_21996_n12996.t3 a_21892_n9816 VSS.t3571 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X557 a_26844_n20485 a_26756_n20388 VSS.t2089 VSS.t2088 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X558 a_27316_n14820 a_21996_n12996.t4 a_26563_n12212 VSS.t3572 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X559 VDD.t1507 a_27744_n12908 a_27639_n12537 VDD.t1506 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X560 VDD.t2110 a_43725_908 a_43845_376 VDD.t2109 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X561 a_40652_n1572 a_40196_n1884 VDD.t1661 VDD.t1660 pfet_06v0 ad=0.5368p pd=3.32u as=0.35315p ps=1.96u w=1.22u l=0.5u
X562 a_11023_n20230.t19 a_13623_n20230.t19 VDD.t578 VDD.t577 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X563 VSS.t3 a_22444_332.t13 a_40859_2428 VSS.t2 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X564 VSS.t1855 a_28456_n364 a_28352_n320 VSS.t1854 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X565 VSS.t2421 a_24236_2258.t3 a_22444_2253.t3 VSS.t2420 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X566 a_34708_n5896.t6 a_33776_n5896.t10 VSS.t874 VSS.t873 nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X567 a_24604_n20485 a_24516_n20388 VSS.t1734 VSS.t1733 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X568 VDD.t1659 a_36388_1944 a_37024_1944.t7 VDD.t1658 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X569 a_30468_n3844 a_27259_804.t3 a_29444_n4328.t0 VSS.t850 nfet_06v0 ad=0.1517p pd=1.19u as=0.2132p ps=1.34u w=0.82u l=0.6u
X570 a_22220_n9860 a_24716_n5156.t3 a_24180_n5112 VSS.t1376 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X571 VSS.t144 a_33496_n6659.t11 a_31628_n5940.t14 VSS.t143 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X572 a_24716_n5156.t0 a_24233_n8684 VSS.t1061 VSS.t1060 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X573 a_27516_n20052 a_27428_n20008 VSS.t3567 VSS.t3566 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X574 VSS.t3981 a_29408_1944.t9 OUT[0].t6 VSS.t3980 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X575 a_27932_n3543 a_28144_n4708 a_28225_n4327 VDD.t3757 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X576 VDD.t2754 a_36588_n9509 a_36500_n9412 VDD.t2753 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X577 a_21692_n20052 a_21604_n20008 VSS.t3518 VSS.t1164 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X578 a_30584_n11296 a_29744_n10980 a_30296_n10980 VSS.t3669 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X579 a_23072_n13432.t3 a_29744_n15604.t10 VSS.t1722 VSS.t1721 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X580 a_29408_1944.t3 a_22052_1944 VSS.t2796 VSS.t2795 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X581 a_40299_n2276 a_28009_n1192.t2 a_26060_n878.t1 VSS.t3556 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X582 a_39500_n12645 a_39412_n12548 VSS.t1965 VSS.t1964 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X583 VDD.t3056 a_38268_n20052 a_38180_n20008 VDD.t3011 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X584 a_24128_n10112 a_22016_n10529 a_23816_n10112 VDD.t1880 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X585 VDD.t1762 a_44092_n16916 a_44004_n16872 VDD.t1761 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X586 VSS.t1724 a_29744_n15604.t11 a_23072_n13432.t2 VSS.t1723 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X587 VDD.t793 a_25612_n878.t2 a_27706_n1572 VDD.t792 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X588 a_11087_n7460.t0 a_13623_n6840.t18 a_13501_n6460.t0 VSS.t721 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X589 a_31548_n10172.t6 a_33496_n8222.t8 VSS.t294 VSS.t293 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X590 a_31656_n704 a_29856_n1121 a_30716_n1148 VSS.t1006 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X591 VDD.t3382 a_44092_n13780 a_44004_n13736 VDD.t3381 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X592 VDD.t3062 a_40196_1944 a_41392_1944.t6 VDD.t3061 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X593 a_30808_n10600 a_30136_n10600 VDD.t1204 VDD.t1203 pfet_06v0 ad=0.3172p pd=1.74u as=0.4005p ps=2.12u w=1.22u l=0.5u
X594 VSS.t411 a_11023_n17552.t23 a_11087_n18172.t28 VSS.t60 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X595 a_29076_n8292.t2 a_25019_n3588.t2 a_33780_n5112 VSS.t3472 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X596 VDD.t3067 a_30036_n7464 a_30740_n7464 VDD.t3066 pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X597 VDD.t286 a_33496_n8222.t9 a_31548_n10172.t15 VDD.t285 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X598 VDD.t3573 a_39724_n11077 a_39636_n10980 VDD.t3572 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X599 a_43728_1248 a_41616_1564 a_43416_1248 VDD.t2747 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X600 a_30408_n1104 a_29444_n708 a_30204_n1104 VSS.t2818 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X601 a_41180_n20485 a_41092_n20388 VSS.t2788 VSS.t2787 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X602 EOC.t6 a_45648_1564.t11 VSS.t31 VSS.t30 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X603 a_40060_n20485 a_39972_n20388 VSS.t3456 VSS.t3455 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X604 a_24220_n15260 a_23912_n15216 VSS.t1005 VSS.t1004 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X605 VDD.t50 a_45648_1564.t12 EOC.t13 VDD.t49 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X606 a_44092_n20052 a_44004_n20008 VSS.t3511 VSS.t3510 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X607 VDD.t1635 a_35356_n18484 a_35268_n18440 VDD.t1634 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X608 a_27485_n10068 a_25573_n12167 VSS.t2172 VSS.t2171 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
D15 a_23072_n13432.t20 VDD.t471 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X609 a_34860_n3189 a_34552_n3140 VSS.t1866 VSS.t1865 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X610 a_11087_n18172.t30 a_2167_3472.t80 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X611 a_37785_n364 a_37368_n320 a_38161_n320 VSS.t1802 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X612 a_47004_n1669 a_46916_n1572 VSS.t2232 VSS.t2231 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X613 VDD.t3022 a_27337_n3140 a_28225_n4327 VDD.t3021 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
D16 VSS.t770 a_24481_761.t19 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X614 VDD.t3944 a_33116_n18484 a_33028_n18440 VDD.t3943 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X615 a_30372_376 a_29812_860 a_30244_860 VSS.t3594 nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X616 VDD.t162 a_33496_n6659.t12 a_31628_n5940.t29 VDD.t161 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X617 VSS.t2751 a_11023_n4162.t21 VSS.t2751 VSS.t66 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.28u
X618 a_23207_n4708 a_23479_n5156 a_23228_n6679 VDD.t2240 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X619 VDD.t2574 a_37372_n5940 a_37284_n5896 VDD.t2573 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X620 a_22016_n1121 a_21604_n708 VSS.t3437 VSS.t3436 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X621 a_31455_n13648 a_30555_n13780 VDD.t1625 VDD.t1624 pfet_06v0 ad=0.1313p pd=1.025u as=0.29465p ps=1.74u w=0.505u l=0.5u
X622 VDD.t1689 a_37024_1944.t9 OUT[2].t14 VDD.t1688 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X623 VDD.t1096 a_22220_n9860 a_22116_n9412 VDD.t1095 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X624 VDD.t3956 a_31235_n9860 a_29992_n11150 VDD.t3955 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X625 a_32628_n10512 a_31460_n10116 a_32424_n10512 VDD.t1279 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X626 VDD.t1589 a_21772_n452.t5 a_13623_n22908.t1 VDD.t1588 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X627 a_40956_n4372 a_40868_n4328 VSS.t2654 VSS.t2653 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X628 a_39500_n7941 a_39412_n7844 VSS.t2941 VSS.t2940 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X629 a_11023_n4162.t8 a_13623_n4162.t17 VSS.t570 VSS.t569 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X630 VDD.t2913 a_47452_n7508 a_47364_n7464 VDD.t2912 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X631 VDD.t3876 a_27180_n18484 a_27092_n18440 VDD.t3875 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X632 a_46220_n17349 a_46132_n17252 VSS.t1262 VSS.t1261 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X633 VSS.t1349 a_13623_n14874.t18 a_11023_n14874.t2 VSS.t1348 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X634 a_10712_4516.t2 a_3935_4156.t5 VSS.t454 VSS.t382 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X635 a_26907_n616 a_26431_n1192 VSS.t3277 VSS.t3276 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X636 VDD.t3748 a_47452_n4372 a_47364_n4328 VDD.t3747 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X637 a_11087_n20850.t2 a_11023_n20230.t22 VSS.t1923 VSS.t62 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X638 a_46220_n14213 a_46132_n14116 VSS.t1215 VSS.t1214 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X639 a_n199_2852 a_n263_3472.t16 VSS.t2084 VSS.t2083 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X640 a_37372_n9076 a_37284_n9032 VSS.t3392 VSS.t3391 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X641 a_42860_n5940 a_42772_n5896 VSS.t3333 VSS.t3332 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X642 a_28435_n10599 a_28519_n10160.t3 a_28455_n10116 VSS.t839 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X643 VSS.t841 a_28519_n10160.t4 a_28721_n9076.t0 VSS.t840 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X644 a_38268_n20485 a_38180_n20388 VSS.t3093 VSS.t3092 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X645 a_11023_n17552.t8 a_13623_n17552.t17 VSS.t77 VSS.t76 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X646 VDD.t427 a_33216_1944.t12 OUT[1].t12 VDD.t426 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X647 VSS.t192 a_11023_n22908.t21 a_11087_n23528.t29 VSS.t64 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X648 a_22464_n7393 a_22052_n6980 VDD.t1491 VDD.t1490 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X649 a_11087_n23528.t31 a_2167_3472.t71 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X650 VSS.t79 a_13623_n17552.t18 a_11023_n17552.t7 VSS.t78 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X651 a_23004_n2332 a_27259_804.t4 VDD.t799 VDD.t798 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X652 VDD.t3354 a_42636_n9509 a_42548_n9412 VDD.t3353 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X653 VSS.t714 a_21772_n20836.t10 a_13623_n6840.t7 VSS.t713 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X654 a_11087_n23528.t28 a_11023_n22908.t22 VSS.t193 VSS.t66 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X655 a_24069_n12398 a_23949_n12996 VDD.t1194 VDD.t1193 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
D17 VSS.t3776 XRST.t0 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X656 VSS.t723 a_13623_n6840.t19 a_11023_n6840.t2 VSS.t722 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X657 a_25817_804 a_24913_864 VDD.t2937 VDD.t2936 pfet_06v0 ad=0.3432p pd=2.44u as=0.3276p ps=1.62u w=0.78u l=0.5u
X658 a_22444_332.t2 a_25836_n1236.t8 VDD.t1071 VDD.t1070 pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X659 VDD.t3699 a_27337_1944.t2 a_22820_n2804 VDD.t3698 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X660 a_32359_n4372 a_33015_n4284 a_32911_n4240 VDD.t2814 pfet_06v0 ad=0.25375p pd=1.51u as=0.1313p ps=1.025u w=0.505u l=0.5u
D18 a_22220_690.t5 VDD.t778 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X661 VSS.t146 a_33496_n6659.t13 a_31628_n5940.t13 VSS.t145 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X662 a_43084_n9509 a_42996_n9412 VSS.t1917 VSS.t1916 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X663 VSS.t1825 a_13623_n12196.t18 a_11023_n12196.t2 VSS.t1824 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X664 a_46668_n18917 a_46580_n18820 VSS.t3037 VSS.t3036 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X665 a_39164_n4805 a_39076_n4708 VSS.t2865 VSS.t2864 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X666 a_27302_n9816 a_26470_n9322 a_27154_n9240 VDD.t996 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X667 VSS.t772 a_24481_761.t20 a_29744_n15604.t2 VSS.t771 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X668 a_11087_n15494.t0 a_13623_n14874.t19 a_13501_n14494.t0 VSS.t1350 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X669 VDD.t1788 a_21692_n15781 a_21604_n15684 VDD.t1787 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X670 VDD.t668 a_13623_n6840.t20 a_11023_n6840.t3 VDD.t667 pfet_03v3 ad=1.82p pd=6.9u as=0.728p ps=3.32u w=2.8u l=0.28u
X671 a_44428_n18917 a_44340_n18820 VSS.t2041 VSS.t2040 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X672 VSS.t308 a_21772_n11428.t8 a_13623_n14874.t7 VSS.t307 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X673 a_13501_n17172.t9 a_13623_n17552.t19 a_11087_n18172.t9 VSS.t80 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X674 VDD.t2582 a_45100_1467 a_45012_1564 VDD.t2581 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X675 VDD.t4237 a_27852_n18917 a_27764_n18820 VDD.t4236 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X676 a_31960_n13648 a_31664_n13292 a_30903_n13780 VDD.t1728 pfet_06v0 ad=0.2424p pd=1.465u as=0.25375p ps=1.51u w=0.505u l=0.5u
X677 a_31799_n7508 a_32560_n7020 a_32351_n7376 VSS.t1331 nfet_06v0 ad=0.2007p pd=1.475u as=94.5f ps=0.885u w=0.36u l=0.6u
X678 a_43532_n7941 a_43444_n7844 VSS.t3265 VSS.t3264 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X679 a_37484_n17349 a_37396_n17252 VSS.t1587 VSS.t1586 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X680 a_32720_n13248 a_23072_n13432.t21 VSS.t488 VSS.t487 nfet_06v0 ad=43.199997f pd=0.6u as=0.2016p ps=1.48u w=0.36u l=0.6u
X681 a_13623_n17552.t5 a_21772_n8292.t10 VSS.t433 VSS.t432 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X682 VDD.t3270 a_28524_n17349 a_28436_n17252 VDD.t3269 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X683 OUT[0].t5 a_29408_1944.t10 VSS.t3983 VSS.t3982 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X684 VDD.t714 a_24481_761.t21 a_39804_464 VDD.t713 pfet_06v0 ad=0.45p pd=2.02u as=0.3432p ps=2.44u w=0.78u l=0.5u
X685 a_27646_n4558 a_27190_n5112 a_27414_n5112 VDD.t1157 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X686 VDD.t1970 a_25612_n18917 a_25524_n18820 VDD.t1969 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X687 a_37484_n14213 a_37396_n14116 VSS.t2509 VSS.t2508 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X688 a_36120_n4 a_35568_n4 a_35916_n4 VDD.t4013 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X689 VDD.t3044 a_40956_n12212 a_40868_n12168 VDD.t3043 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X690 VSS.t296 a_33496_n8222.t10 a_31548_n10172.t5 VSS.t295 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X691 a_28225_n9031 a_25972_n6276 a_28617_n8548 VDD.t1795 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X692 VDD.t3950 a_43084_n11077 a_42996_n10980 VDD.t3949 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X693 a_35244_n17349 a_35156_n17252 VSS.t957 VSS.t956 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X694 a_32560_n7020 a_31548_n10172.t16 VSS.t282 VSS.t281 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X695 a_35244_n14213 a_35156_n14116 VSS.t1492 VSS.t1491 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X696 EOC.t12 a_45648_1564.t13 VDD.t52 VDD.t51 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X697 VDD.t2783 a_43420_n2804 a_43332_n2760 VDD.t2782 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X698 a_44540_n7508 a_44452_n7464 VSS.t2968 VSS.t2967 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X699 VDD.t2617 a_21692_n13308.t16 a_21940_n11684 VDD.t2616 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X700 a_11087_n20850.t31 a_2167_3472.t17 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X701 a_34188_n5112 a_25019_n3588.t3 a_29076_n8292.t2 VSS.t3473 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X702 a_11023_n9518.t18 a_13623_n9518.t12 VDD.t256 VDD.t255 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X703 VDD.t3088 a_38716_n10644 a_38628_n10600 VDD.t3087 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X704 a_47452_n12212 a_47364_n12168 VSS.t1180 VSS.t1179 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X705 a_11087_n12816.t20 a_13623_n12196.t19 a_13501_n11816.t10 VSS.t1826 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X706 a_22588_n15781 a_22500_n15684 VSS.t3023 VSS.t3022 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X707 VDD.t552 a_13623_n4162.t18 a_11023_n4162.t19 VDD.t551 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X708 a_34344_n3840 a_33416_n4240 a_34176_n3840 VSS.t3169 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X709 OUT[4].t15 a_41392_1944.t8 VDD.t1373 VDD.t1372 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X710 VSS.t2673 a_21692_n13308.t17 a_22052_n6980 VSS.t2672 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X711 a_27792_n320 a_24481_761.t22 VSS.t774 VSS.t773 nfet_06v0 ad=43.199997f pd=0.6u as=0.2016p ps=1.48u w=0.36u l=0.6u
X712 a_47452_n1669 a_47364_n1572 VSS.t1142 VSS.t1141 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D19 VSS.t335 a_10712_4516.t31 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X713 a_45212_n12212 a_45124_n12168 VSS.t3025 VSS.t3024 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X714 VDD.t2045 a_39612_n20052 a_39524_n20008 VDD.t2044 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D20 a_23072_n13432.t22 VDD.t472 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X715 a_22116_860 a_22444_332.t14 a_22096_376 VSS.t4 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X716 a_31076_376 a_30372_376 VSS.t4015 VSS.t4014 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X717 a_31376_n6592 a_23072_n13432.t23 VSS.t490 VSS.t489 nfet_06v0 ad=43.199997f pd=0.6u as=0.2016p ps=1.48u w=0.36u l=0.6u
X718 a_32424_n10512 a_31872_n10529 a_32220_n10512 VDD.t3750 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X719 VSS.t3296 a_26239_n12996 a_26175_n12951 VSS.t3295 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X720 VDD.t2943 a_42300_n7508 a_42212_n7464 VDD.t2942 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X721 VSS.t33 a_45648_1564.t14 EOC.t5 VSS.t32 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X722 VDD.t2072 a_42300_n4372 a_42212_n4328 VDD.t2071 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X723 a_27302_n9816 a_26470_n9322 a_27134_n9816 VSS.t3214 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X724 VDD.t2865 a_48012_n18917 a_47924_n18820 VDD.t2864 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X725 a_38716_n16916 a_38628_n16872 VSS.t2964 VSS.t2963 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X726 a_22772_n1104 a_21604_n708 a_22568_n1104 VDD.t3360 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X727 a_34840_n3456 a_34000_n3140 a_34552_n3140 VSS.t2776 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X728 a_22772_n8944 a_23072_n13432.t24 VDD.t474 VDD.t473 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X729 a_31760_n12168 a_30787_n12167 VDD.t1835 VDD.t1834 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X730 a_31772_n16916 a_31684_n16872 VSS.t2960 VSS.t2959 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X731 a_23728_464 a_23136_447 a_23524_464 VDD.t1895 pfet_06v0 ad=0.19315p pd=1.27u as=0.1313p ps=1.025u w=0.505u l=0.5u
X732 a_22772_n5808 a_23072_n13432.t25 VDD.t476 VDD.t475 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X733 VDD.t2492 a_37820_n18484 a_37732_n18440 VDD.t2491 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X734 VSS.t1726 a_29744_n15604.t12 a_23072_n13432.t4 VSS.t1725 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X735 a_13501_n19850.t18 a_13623_n20230.t20 a_11087_n20850.t28 VSS.t618 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X736 a_13501_n22528.t18 a_11023_n22908.t23 a_11087_n23528.t12 VDD.t207 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X737 VDD.t1766 a_28456_n364 a_28352_n320 VDD.t1765 pfet_06v0 ad=0.3432p pd=2.44u as=0.2028p ps=1.3u w=0.78u l=0.5u
X738 a_28225_n9031 a_24492_n5156 VDD.t3497 VDD.t415 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X739 VDD.t1673 a_28009_n12168 a_29360_n12864 VDD.t1672 pfet_06v0 ad=0.3432p pd=2.44u as=0.2028p ps=1.3u w=0.78u l=0.5u
D21 XRST.t1 VDD.t3700 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X740 VDD.t2895 a_36700_n18484 a_36612_n18440 VDD.t2894 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X741 VSS.t1209 a_25237_n4327 a_25759_n3544 VSS.t1208 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X742 a_13501_n6460.t1 a_13623_n6840.t21 a_11087_n7460.t1 VSS.t724 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X743 VSS.t4268 a_28568_n16066 a_23564_n17700 VSS.t4267 nfet_06v0 ad=0.151p pd=1.185u as=0.1261p ps=1.005u w=0.485u l=0.6u
X744 a_36388_n1572 a_35940_n1931 VSS.t3111 VSS.t3110 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X745 a_40260_n408 a_39556_n4 VDD.t3288 VDD.t3287 pfet_06v0 ad=0.3477p pd=1.79u as=0.4392p ps=1.94u w=1.22u l=0.5u
X746 a_27531_n11593 a_27055_n12168 a_27279_n12146 VSS.t2918 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X747 a_13501_n22528.t8 a_13623_n22908.t12 a_11087_n23528.t8 VSS.t207 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X748 a_42748_n18484 a_42660_n18440 VSS.t2958 VSS.t2957 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X749 a_23220_n7376 a_23072_n13432.t26 VDD.t478 VDD.t477 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X750 a_42748_n15348 a_42660_n15304 VSS.t3418 VSS.t3417 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X751 a_23004_n2332 a_25836_n1236.t9 VDD.t1073 VDD.t1072 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X752 a_40508_n18484 a_40420_n18440 VSS.t2494 VSS.t2493 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X753 a_29744_n15604.t6 a_24481_761.t23 VDD.t716 VDD.t715 pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X754 a_13623_n20230.t14 a_21772_n3588.t6 VDD.t574 VDD.t573 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X755 VDD.t1176 a_23564_n8292 a_21772_n8292.t6 VDD.t1175 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X756 a_40508_n15348 a_40420_n15304 VSS.t2935 VSS.t2934 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X757 a_n199_2852 VIN.t0 a_137_4292 VSS.t3091 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X758 VDD.t1685 a_43644_n15348 a_43556_n15304 VDD.t1684 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X759 a_42412_n101 a_42324_n4 VSS.t3416 VSS.t3415 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X760 a_22364_n1104 a_22264_n1148.t2 VDD.t3711 VDD.t3710 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
D22 a_23072_n13432.t27 VDD.t479 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X761 a_41628_n2804 a_41540_n2760 VSS.t3384 VSS.t3383 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X762 VDD.t3962 a_29211_n6724 a_29123_n6679 VDD.t3961 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X763 VDD.t3099 a_44428_n6373 a_44340_n6276 VDD.t3098 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X764 a_32712_n10112 a_31872_n10529 a_32424_n10512 VSS.t3823 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X765 VDD.t3321 a_44428_n3237 a_44340_n3140 VDD.t3320 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X766 a_25600_n5895 a_21692_n6694.t9 a_25620_n5412 VSS.t679 nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X767 a_22568_n10512 a_22016_n10529 a_22364_n10512 VDD.t1879 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X768 a_35356_n12212 a_35268_n12168 VSS.t3240 VSS.t3239 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X769 VDD.t2901 a_41404_n15348 a_41316_n15304 VDD.t2900 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D23 a_24481_761.t24 VDD.t717 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X770 VSS.t2752 a_11023_n4162.t22 VSS.t2752 VSS.t68 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.28u
X771 VDD.t4155 a_34652_n11391 a_34538_n10980 VDD.t4154 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X772 VDD.t3161 a_39276_n18917 a_39188_n18820 VDD.t3160 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X773 VDD.t3387 a_27516_n20052 a_27428_n20008 VDD.t3386 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X774 VDD.t3267 a_34460_n16916 a_34372_n16872 VDD.t3266 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X775 VDD.t88 a_13623_n17552.t20 a_11023_n17552.t19 VDD.t87 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X776 a_23319_n2759 a_22500_n1976 a_23507_n2759 VDD.t1702 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X777 a_31628_n5940.t12 a_33496_n6659.t14 VSS.t148 VSS.t147 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
D24 a_23072_n13432.t28 VDD.t480 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X778 VDD.t3775 a_21692_n20052 a_21604_n20008 VDD.t3774 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X779 a_39612_n20485 a_39524_n20388 VSS.t3379 VSS.t3378 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X780 a_23036_n18917 a_22948_n18820 VSS.t3425 VSS.t3012 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X781 a_35692_n15348 a_35604_n15304 VSS.t2249 VSS.t2248 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X782 a_31965_n8292 a_29123_n6679 VSS.t2603 VSS.t2602 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X783 a_27123_n12872 a_26983_n12728 a_26635_n12996 VSS.t3969 nfet_06v0 ad=0.134p pd=1.1u as=0.176p ps=1.68u w=0.4u l=0.6u
X784 VDD.t2812 a_37036_n18917 a_36948_n18820 VDD.t2811 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X785 VSS.t2891 a_25577_n14956 a_25472_n14816 VSS.t2890 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X786 VDD.t1657 a_36388_1944 a_37024_1944.t6 VDD.t1656 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X787 a_43980_n7941 a_43892_n7844 VSS.t1931 VSS.t1930 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X788 VDD.t3241 a_32220_n16916 a_32132_n16872 VDD.t3240 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X789 VDD.t4047 a_25685_n7463 a_26095_n7464 VDD.t4046 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X790 VDD.t956 a_27485_n8500 a_27605_n9032 VDD.t955 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X791 a_33452_n15348 a_33364_n15304 VSS.t2929 VSS.t2831 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X792 a_35244_n13780 a_35156_n13736 VSS.t3345 VSS.t3344 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X793 a_27055_n12168 a_26431_n12168 a_26907_n11592 VSS.t3261 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X794 VSS.t2539 a_27302_n13160 a_27778_n13161 VSS.t2538 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X795 VSS.t931 a_32636_n2020 a_32100_n1976 VSS.t930 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X796 VDD.t3170 a_30092_n18917 a_30004_n18820 VDD.t3169 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X797 VSS.t3050 a_34428_n452.t2 a_34380_n408 VSS.t3049 nfet_06v0 ad=0.2132p pd=1.34u as=98.399994f ps=1.06u w=0.82u l=0.6u
X798 VDD.t482 a_23072_n13432.t29 a_31068_n6276 VDD.t481 pfet_06v0 ad=0.45p pd=2.02u as=0.3432p ps=2.44u w=0.78u l=0.5u
X799 VDD.t1742 a_13623_n12196.t20 a_11023_n12196.t3 VDD.t1741 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X800 VDD.t444 a_34708_n5896.t16 a_33496_n8222.t6 VDD.t443 pfet_06v0 ad=0.3608p pd=2.52u as=0.2952p ps=1.54u w=0.82u l=0.5u
X801 a_29408_1944.t2 a_22052_1944 VSS.t2794 VSS.t2793 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X802 VSS.t999 a_39648_n2020 a_23564_1116.t0 VSS.t998 nfet_06v0 ad=0.2344p pd=1.56u as=0.3608p ps=2.52u w=0.82u l=0.6u
X803 a_25057_n6976 a_23072_n13432.t30 VSS.t492 VSS.t491 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X804 a_32220_n10512 a_30808_n10116 VDD.t2867 VDD.t2866 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X805 a_11023_n12196.t4 a_13623_n12196.t21 VDD.t1744 VDD.t1743 pfet_03v3 ad=0.728p pd=3.32u as=1.82p ps=6.9u w=2.8u l=0.28u
X806 a_34460_n20052 a_34372_n20008 VSS.t3409 VSS.t3408 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X807 VDD.t2175 a_25724_n18484 a_25636_n18440 VDD.t2174 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X808 VSS.t2949 a_35848_n3868 a_23564_n3588.t0 VSS.t2948 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X809 VSS.t1878 a_25972_n6276 a_28841_n8548 VSS.t1877 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X810 VDD.t2254 a_43196_n10644 a_43108_n10600 VDD.t2253 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X811 VDD.t484 a_23072_n13432.t31 a_28492_n12548 VDD.t483 pfet_06v0 ad=0.45p pd=2.02u as=0.3432p ps=2.44u w=0.78u l=0.5u
X812 a_32780_n2672 a_31392_n2760 VSS.t4219 VSS.t4218 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X813 VSS.t4318 a_26266_n13736 a_26742_n13160 VSS.t4317 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X814 VDD.t3851 a_22876_n13692 a_22772_n13648 VDD.t3850 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X815 VSS.t1015 a_27485_n8500 a_27605_n8456 VSS.t1014 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X816 VSS.t4134 a_22140_n6694.t4 a_25020_n11383 VSS.t4133 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X817 a_32220_n20052 a_32132_n20008 VSS.t3403 VSS.t3402 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X818 VSS.t610 a_21772_n3588.t7 a_13623_n20230.t6 VSS.t609 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X819 VDD.t3263 a_39276_n9509 a_39188_n9412 VDD.t3262 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X820 VDD.t1302 a_13623_n14874.t20 a_11023_n14874.t3 VDD.t1301 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X821 a_23004_n2332 a_27259_804.t5 a_27175_860 VSS.t851 nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X822 a_28040_n12493 a_27639_n12537 a_26983_n12728 VSS.t2156 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X823 VDD.t901 a_44092_n20052 a_44004_n20008 VDD.t900 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X824 a_22876_n13692 a_22568_n13648 VDD.t3792 VDD.t3791 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X825 a_34576_1204 a_32108_n2332.t16 VDD.t4124 VDD.t4123 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X826 a_34068_n4 a_29900_760.t5 a_33920_n4 VDD.t3033 pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X827 a_39612_n4372 a_39524_n4328 VSS.t4072 VSS.t4071 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X828 a_26060_n878.t0 a_28009_n1192.t3 VDD.t3472 VDD.t3471 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X829 VDD.t1886 a_26154_n4536 a_26590_n4536 VDD.t1885 pfet_06v0 ad=0.1656p pd=1.28u as=61.199993f ps=0.7u w=0.36u l=0.5u
X830 a_25975_n184 a_26736_n364 a_26527_51 VSS.t1528 nfet_06v0 ad=0.2007p pd=1.475u as=94.5f ps=0.885u w=0.36u l=0.6u
X831 a_26488_1564 a_25936_1564 a_26284_1564 VDD.t1428 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X832 VDD.t54 a_45648_1564.t15 EOC.t11 VDD.t53 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X833 a_33831_n1400 a_33375_n1976 VDD.t1955 VDD.t1954 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X834 VSS.t3837 a_25237_n5895 a_25530_n5112 VSS.t3836 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X835 a_29360_n12864 a_27639_n12537 a_28232_n12606 VDD.t2083 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X836 a_43196_n16916 a_43108_n16872 VSS.t3019 VSS.t3018 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X837 VSS.t1595 a_31787_n3969 a_29920_n3900.t0 VSS.t1594 nfet_06v0 ad=0.3586p pd=2.51u as=0.2119p ps=1.335u w=0.815u l=0.6u
X838 a_25940_n17606.t0 a_32262_n452 VSS.t1446 VSS.t1445 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
D25 a_23072_n13432.t32 VDD.t485 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X839 VDD.t1375 a_41392_1944.t9 OUT[4].t14 VDD.t1374 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X840 VSS.t2665 a_26328_n6654.t12 a_21692_n13308.t5 VSS.t2664 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X841 VDD.t3754 a_29540_n11728 a_24492_n5156 VDD.t3753 pfet_06v0 ad=0.389p pd=2.02u as=0.5368p ps=3.32u w=1.22u l=0.5u
X842 VDD.t2832 a_47004_n18484 a_46916_n18440 VDD.t2831 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X843 VSS.t853 a_27259_804.t6 a_27628_n3841 VSS.t852 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X844 VSS.t2559 a_35392_n10172 a_28519_n10160.t0 VSS.t2558 nfet_06v0 ad=0.2344p pd=1.56u as=0.3608p ps=2.52u w=0.82u l=0.6u
X845 a_29756_n20485 a_29668_n20388 VSS.t2850 VSS.t2849 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X846 VDD.t4269 a_23484_n16916 a_23396_n16872 VDD.t4268 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X847 VSS.t1188 a_25237_n13735 a_25642_n13736 VSS.t1187 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X848 a_27511_n1170 a_27055_n1192 a_27279_n1170 VDD.t3116 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X849 VDD.t1154 a_36217_n3500 a_36112_n3456 VDD.t1153 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X850 a_27259_804.t0 a_30452_n5156.t4 VSS.t1078 VSS.t1077 nfet_06v0 ad=0.2255p pd=1.37u as=0.3608p ps=2.52u w=0.82u l=0.6u
X851 a_30320_n6636 a_31548_n10172.t17 VDD.t276 VDD.t275 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X852 a_11023_n22908.t18 a_13623_n22908.t13 VDD.t219 VDD.t218 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X853 VDD.t2834 a_40060_n18484 a_39972_n18440 VDD.t2833 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X854 a_26742_n9816 a_26266_n9240 a_26470_n9322 VSS.t3542 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X855 a_22444_2253.t6 a_24236_2258.t4 VDD.t2335 VDD.t2334 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X856 a_42636_n4805 a_42548_n4708 VSS.t2327 VSS.t2326 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X857 a_28121_n10980 a_27391_n11384 VDD.t3596 VDD.t3595 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X858 VSS.t3197 a_35288_n1975 a_34248_n3310 VSS.t3196 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X859 a_36709_n2276 a_34953_n1572 VSS.t2881 VSS.t2880 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X860 a_22364_n10512 a_22264_n10556 VDD.t2177 VDD.t2176 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X861 a_11087_n23528.t32 a_2167_3472.t70 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X862 VDD.t1917 a_27281_n16854 a_29180_n9387 VDD.t1916 pfet_06v0 ad=0.5913p pd=3.27u as=0.2847p ps=1.615u w=1.095u l=0.5u
X863 a_23484_n20052 a_23396_n20008 VSS.t3313 VSS.t2556 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X864 VDD.t3157 a_44876_n15781 a_44788_n15684 VDD.t3156 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X865 VDD.t3002 a_44876_n6373 a_44788_n6276 VDD.t3001 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X866 VDD.t429 a_33216_1944.t13 OUT[1].t11 VDD.t428 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X867 VDD.t2941 a_44876_n12645 a_44788_n12548 VDD.t2940 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X868 a_27758_n13714 a_27302_n13160 a_27526_n13714 VDD.t2461 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X869 VDD.t2308 a_44876_n3237 a_44788_n3140 VDD.t2307 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X870 a_43644_n4372 a_43556_n4328 VSS.t3958 VSS.t3957 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X871 a_37680_n320 a_35156_n325 a_37368_n320 VSS.t3066 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X872 VDD.t42 a_28156_n6412.t17 a_26440_n5940.t0 VDD.t41 pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X873 a_30092_n10980 a_29992_n11150 VSS.t3027 VSS.t3026 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X874 VDD.t2955 a_42636_n15781 a_42548_n15684 VDD.t2954 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X875 a_32108_n2332.t4 a_35456_n4628.t10 VSS.t4163 VSS.t4162 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X876 VDD.t1536 a_42636_n12645 a_42548_n12548 VDD.t1535 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X877 a_11087_n10138.t3 a_11023_n9518.t23 a_13501_n9138.t2 VDD.t543 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X878 a_28972_n17349 a_28884_n17252 VSS.t1090 VSS.t1089 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X879 VDD.t3368 a_38268_n18484 a_38180_n18440 VDD.t3367 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X880 VDD.t4041 a_45324_n9509 a_45236_n9412 VDD.t4040 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X881 a_22772_n13648 a_21604_n13252 a_22568_n13648 VDD.t2141 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X882 VSS.t2629 a_24573_n6724 a_24693_n6680 VSS.t2628 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
D26 VSS.t493 a_23072_n13432.t33 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X883 a_11023_n20230.t18 a_13623_n20230.t21 VDD.t580 VDD.t579 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X884 OUT[0].t4 a_29408_1944.t11 VSS.t3985 VSS.t3984 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X885 a_11087_n20850.t3 a_11023_n20230.t23 a_13501_n19850.t8 VDD.t1843 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X886 VDD.t2337 a_22444_2253.t9 a_n263_3472.t14 VDD.t453 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X887 a_21692_n5468.t13 a_26440_n5940.t7 VDD.t391 VDD.t390 pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X888 a_37820_n12212 a_37732_n12168 VSS.t2852 VSS.t2851 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X889 a_24569_n11820 a_23072_n13432.t34 VDD.t487 VDD.t486 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X890 a_11087_n7460.t27 a_11023_n6840.t23 a_13501_n6460.t8 VDD.t109 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X891 a_36700_n12212 a_36612_n12168 VSS.t2103 VSS.t2102 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X892 OUT[2].t13 a_37024_1944.t10 VDD.t1691 VDD.t1690 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X893 a_30428_n12645 a_30340_n12548 VSS.t3443 VSS.t3442 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X894 a_28232_n12606 a_27744_n12908 a_28492_n12548 VDD.t1505 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X895 VDD.t3765 a_41068_n5940 a_40980_n5896 VDD.t3764 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X896 VSS.t1643 a_34576_1204 a_34471_1575 VSS.t1642 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X897 a_35371_n617 a_34895_n1192 a_35119_n1170 VSS.t1451 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X898 a_24836_n4708 a_24716_n5156.t4 a_22220_n9860 VDD.t1325 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X899 a_48012_n17349 a_47924_n17252 VSS.t3487 VSS.t3486 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X900 a_46220_n7941 a_46132_n7844 VSS.t3143 VSS.t3142 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X901 a_35595_n8548 a_29900_n10600.t2 a_28852_n8292.t1 VSS.t3944 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
D27 a_24481_761.t25 VDD.t718 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X902 a_48012_n14213 a_47924_n14116 VSS.t3126 VSS.t3125 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X903 a_11087_n15494.t28 a_11023_n14874.t22 VSS.t57 VSS.t56 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X904 a_23507_n2759 a_22500_n1976 a_23527_n2276 VSS.t1792 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X905 VSS.t337 a_10712_4516.t32 a_10778_2852.t0 VSS.t336 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X906 a_44092_n9076 a_44004_n9032 VSS.t3086 VSS.t3085 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X907 VDD.t3894 a_45660_n10644 a_45572_n10600 VDD.t3893 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X908 a_11087_n23528.t33 a_2167_3472.t69 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X909 VDD.t1591 a_21772_n452.t6 a_13623_n22908.t2 VDD.t1590 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X910 VDD.t4039 a_44540_n10644 a_44452_n10600 VDD.t4038 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X911 VSS.t946 a_23564_n20836 a_21772_n20836.t3 VSS.t945 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X912 a_29744_n15604.t5 a_24481_761.t26 VDD.t720 VDD.t719 pfet_06v0 ad=0.2952p pd=1.54u as=0.3608p ps=2.52u w=0.82u l=0.5u
X913 a_43845_952 a_43725_908 a_43101_841 VSS.t2188 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X914 a_11087_n18172.t27 a_11023_n17552.t24 VSS.t412 VSS.t62 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X915 VSS.t1898 CLK.t3 a_33496_n6659.t0 VSS.t1897 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X916 a_11087_n10138.t25 a_13623_n9518.t13 a_13501_n9138.t18 VSS.t244 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X917 a_13623_n6840.t6 a_21772_n20836.t11 VSS.t716 VSS.t715 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X918 a_27281_n16854 a_22140_n6694.t5 a_27301_n16388 VSS.t4135 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X919 VDD.t3055 a_33533_908 a_33653_376 VDD.t3054 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X920 VDD.t2861 a_42300_n10644 a_42212_n10600 VDD.t2860 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X921 a_26692_1564 a_24481_761.t27 VDD.t722 VDD.t721 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X922 VSS.t3790 a_24088_n16087 a_23564_n20836 VSS.t3789 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X923 a_31676_n3544 a_29920_n3900.t8 a_29560_n3544 VSS.t652 nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X924 a_25132_n16432 a_24964_n14116 a_25559_n12548 VDD.t1838 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X925 a_45660_n16916 a_45572_n16872 VSS.t3119 VSS.t3118 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X926 VDD.t2613 a_26328_n6654.t13 a_21692_n13308.t12 VDD.t2612 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X927 a_44540_n16916 a_44452_n16872 VSS.t3335 VSS.t3334 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X928 a_11023_n9518.t17 a_13623_n9518.t14 VDD.t258 VDD.t257 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X929 a_28744_n14432 a_26944_n14116 a_27804_n14165 VSS.t4000 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X930 a_11087_n12816.t8 a_11023_n12196.t22 VSS.t117 VSS.t56 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X931 VSS.t2802 a_25076_n4.t2 a_22892_n5156.t2 VSS.t2801 nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
X932 a_42300_n16916 a_42212_n16872 VSS.t3339 VSS.t3338 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X933 a_41203_n799 a_41533_n727 a_41653_n1170 VDD.t3546 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X934 VDD.t44 a_28156_n6412.t18 a_26440_n5940.t1 VDD.t43 pfet_06v0 ad=0.3608p pd=2.52u as=0.2952p ps=1.54u w=0.82u l=0.5u
X935 VSS.t1754 a_23564_n11428 a_21772_n11428.t3 VSS.t1753 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X936 VDD.t3147 a_29644_n18917 a_29556_n18820 VDD.t3146 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X937 a_13623_n14874.t6 a_21772_n11428.t9 VSS.t310 VSS.t309 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X938 a_28454_n2424 a_28940_n2406.t2 VDD.t3721 VDD.t3720 pfet_06v0 ad=0.5368p pd=3.32u as=0.4941p ps=2.03u w=1.22u l=0.5u
X939 a_39276_n17349 a_39188_n17252 VSS.t2828 VSS.t2827 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X940 VSS.t395 a_21692_n5468.t18 a_21604_n3844 VSS.t394 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X941 a_30240_n7464 a_29476_n6980 a_30036_n7464 VDD.t2268 pfet_06v0 ad=0.4758p pd=2u as=0.3172p ps=1.74u w=1.22u l=0.5u
X942 a_39276_n14213 a_39188_n14116 VSS.t3616 VSS.t3615 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X943 VSS.t776 a_24481_761.t28 a_36576_n320 VSS.t775 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X944 a_34232_n2272 a_32020_n2276 a_33292_n2716 VDD.t2786 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X945 VDD.t3302 a_27404_n18917 a_27316_n18820 VDD.t3301 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X946 VDD.t3989 a_42748_n12212 a_42660_n12168 VDD.t3988 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X947 a_37036_n17349 a_36948_n17252 VSS.t4045 VSS.t4044 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X948 a_42860_n101 a_42772_n4 VSS.t3681 VSS.t3680 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X949 a_28336_376 a_27572_860 a_28132_376 VDD.t1776 pfet_06v0 ad=0.4758p pd=2u as=0.3172p ps=1.74u w=1.22u l=0.5u
X950 a_38435_864 a_38295_332 a_37947_332 VSS.t1228 nfet_06v0 ad=0.134p pd=1.1u as=0.176p ps=1.68u w=0.4u l=0.6u
X951 VDD.t3568 a_45772_n9509 a_45684_n9412 VDD.t3567 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X952 a_37036_n14213 a_36948_n14116 VSS.t2121 VSS.t2120 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X953 a_32351_n7376 a_31451_n7508 VDD.t4174 VDD.t4173 pfet_06v0 ad=0.1313p pd=1.025u as=0.29465p ps=1.74u w=0.505u l=0.5u
X954 VDD.t2708 a_40508_n12212 a_40420_n12168 VDD.t2707 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X955 VDD.t2261 a_46243_769 a_42604_n2020 VDD.t2260 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X956 a_11087_n15494.t18 a_11023_n14874.t23 a_13501_n14494.t18 VDD.t74 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X957 a_29559_n6456 a_30215_n6265 a_30111_n6221 VDD.t1807 pfet_06v0 ad=0.25375p pd=1.51u as=0.1313p ps=1.025u w=0.505u l=0.5u
X958 VSS.t1341 a_30396_n7508 a_30348_n6980 VSS.t1340 nfet_06v0 ad=0.2132p pd=1.34u as=98.399994f ps=1.06u w=0.82u l=0.6u
X959 a_25577_n14956 a_23072_n13432.t35 VDD.t489 VDD.t488 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X960 a_13501_n6460.t2 a_13623_n6840.t22 a_11087_n7460.t2 VSS.t725 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X961 a_40060_n7508 a_39972_n7464 VSS.t4238 VSS.t4237 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X962 a_34475_n1976 a_33999_n1400 a_34223_n1976 VSS.t3529 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X963 a_22772_n8944 a_21604_n8548 a_22568_n8944 VDD.t3954 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X964 a_47004_n12212 a_46916_n12168 VSS.t3154 VSS.t3153 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X965 a_13501_n17172.t17 a_11023_n17552.t25 a_11087_n18172.t17 VDD.t402 pfet_03v3 ad=1.82p pd=6.9u as=0.728p ps=3.32u w=2.8u l=0.28u
X966 a_44316_n2804 a_44228_n2760 VSS.t3821 VSS.t3504 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X967 a_22016_n6276 a_21916_n6694.t2 a_21812_n6276 VDD.t3494 pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X968 VDD.t3247 a_47116_n6373 a_47028_n6276 VDD.t3246 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X969 a_22772_n5808 a_21604_n5412 a_22568_n5808 VDD.t3496 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X970 a_11087_n20850.t30 a_2167_3472.t14 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X971 VSS.t194 a_11023_n22908.t24 a_11087_n23528.t27 VSS.t68 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X972 a_27700_n14116 a_23072_n13432.t36 VDD.t491 VDD.t490 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X973 VDD.t3046 a_47116_n3237 a_47028_n3140 VDD.t3045 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X974 VDD.t1520 a_34089_n10252 a_33984_n10112 VDD.t1519 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X975 a_40060_n12212 a_39972_n12168 VSS.t4302 VSS.t4301 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X976 VDD.t2219 a_34460_n20052 a_34372_n20008 VDD.t2218 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X977 a_24481_761.t2 a_30192_n15304.t9 VDD.t2284 VDD.t1646 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X978 a_31664_n13292 a_31548_n10172.t18 VSS.t284 VSS.t283 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X979 VDD.t3326 a_32220_n20052 a_32132_n20008 VDD.t3325 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X980 VSS.t1935 a_34068_n4 a_34403_332 VSS.t1934 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X981 a_33564_n16916 a_33476_n16872 VSS.t2329 VSS.t2328 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X982 a_35008_n3456 a_34860_n3189 a_34840_n3456 VSS.t2606 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X983 VDD.t2967 a_39612_n18484 a_39524_n18440 VDD.t2966 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X984 VDD.t3276 a_26172_n14564.t2 a_24965_n9860 VDD.t3275 pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X985 VDD.t4126 a_32108_n2332.t17 a_41204_1243 VDD.t4125 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X986 a_25836_n1236.t3 a_34649_n2412 VSS.t3709 VSS.t3708 nfet_06v0 ad=0.2119p pd=1.335u as=0.3586p ps=2.51u w=0.815u l=0.6u
X987 VSS.t1543 a_29295_n1400 a_29771_n1976 VSS.t1542 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X988 a_29560_n3544 a_29920_n3900.t9 a_32104_n3544 VSS.t653 nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X989 a_24815_n3588.t2 a_29920_n3900.t10 VDD.t600 VDD.t599 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X990 a_11087_n12816.t18 a_11023_n12196.t23 a_13501_n11816.t8 VDD.t128 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X991 a_31324_n16916 a_31236_n16872 VSS.t3176 VSS.t3175 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X992 a_13501_n14494.t1 a_13623_n14874.t21 a_11087_n15494.t1 VSS.t1351 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X993 VDD.t871 a_40652_n1572 a_45648_1564.t6 VDD.t870 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
D28 VSS.t832 a_22220_690.t6 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X994 a_33496_n6659.t2 CLK.t4 VDD.t1817 VDD.t1816 pfet_06v0 ad=0.2542p pd=1.44u as=0.428p ps=2.02u w=0.82u l=0.5u
X995 a_11087_n15494.t2 a_13623_n14874.t22 a_13501_n14494.t2 VSS.t1352 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X996 a_32413_n14564 a_28752_n15348 VDD.t3128 VDD.t3127 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X997 VSS.t1275 a_25612_n6679 a_25524_n6635 VSS.t1274 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X998 a_24609_n8544 a_23072_n13432.t37 VSS.t495 VSS.t494 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X999 VDD.t801 a_27259_804.t7 a_22444_332.t3 VDD.t800 pfet_06v0 ad=0.30535p pd=1.605u as=0.52205p ps=2.045u w=0.985u l=0.5u
X1000 a_11087_n23528.t34 a_2167_3472.t68 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X1001 a_24609_n5408 a_23072_n13432.t38 VSS.t497 VSS.t496 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X1002 a_29659_n14820 a_28121_n10980 a_27852_n14990 VSS.t3685 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1003 a_31685_n9262 a_31565_n9860 VDD.t2213 VDD.t2212 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X1004 a_13501_n17172.t8 a_13623_n17552.t21 a_11087_n18172.t8 VSS.t81 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1005 a_40652_n1572 a_40196_n1884 VSS.t1744 VSS.t1743 nfet_06v0 ad=0.3608p pd=2.52u as=0.2344p ps=1.56u w=0.82u l=0.6u
X1006 a_22364_n8944 a_22264_n8988 VDD.t2923 VDD.t2922 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X1007 a_22364_n5808 a_22264_n5852 VDD.t1526 VDD.t1525 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X1008 a_29744_n10980 a_29332_n11301 VSS.t3559 VSS.t3558 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1009 VDD.t2903 a_46556_n15348 a_46468_n15304 VDD.t2902 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1010 a_10778_2852.t1 a_10712_4516.t33 VDD.t326 VDD.t325 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1011 VDD.t1377 a_41392_1944.t10 OUT[4].t13 VDD.t1376 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1012 a_23703_n5156.t1 a_28454_n2424 VDD.t3257 VDD.t3256 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1013 VDD.t1841 a_41740_n7941 a_41652_n7844 VDD.t1840 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1014 a_24573_n9860 a_24965_n9860 VDD.t1981 VDD.t996 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1015 a_38268_n12212 a_38180_n12168 VSS.t2149 VSS.t2148 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1016 a_39352_464 a_38951_420 a_38295_332 VSS.t3300 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1017 a_2167_3472.t0 a_13623_n4162.t19 VSS.t572 VSS.t571 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1018 VSS.t3687 a_25880_n11708 a_21692_n5111.t0 VSS.t3686 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X1019 VDD.t2935 a_41740_n4805 a_41652_n4708 VDD.t2934 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D29 VSS.t4136 a_22140_n6694.t6 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1020 a_13501_n11816.t11 a_13623_n12196.t22 a_11087_n12816.t21 VSS.t1827 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1021 a_27988_n20388 a_27540_n20747 VSS.t2944 VSS.t2943 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X1022 VDD.t1809 a_37585_n3140 a_29263_n3588.t0 VDD.t1808 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1023 a_36588_n9509 a_36500_n9412 VSS.t3671 VSS.t3670 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1024 VDD.t2873 a_37372_n16916 a_37284_n16872 VDD.t2872 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1025 a_13501_n6460.t11 a_11023_n6840.t24 a_11087_n7460.t26 VDD.t110 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1026 a_27623_n10830 a_27167_n10808 a_27391_n11384 VDD.t3569 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X1027 a_11087_n12816.t22 a_13623_n12196.t23 a_13501_n11816.t12 VSS.t1828 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X1028 a_22812_n7376 a_22712_n7420 VDD.t911 VDD.t910 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X1029 a_32220_n10512 a_30808_n10116 VSS.t2931 VSS.t2930 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1030 VDD.t3159 a_36252_n16916 a_36164_n16872 VDD.t3158 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1031 VDD.t3137 a_37372_n13780 a_37284_n13736 VDD.t3136 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1032 a_40508_n9076 a_40420_n9032 VSS.t3731 VSS.t3730 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1033 a_44876_n11077 a_44788_n10980 VSS.t3254 VSS.t3253 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1034 a_28800_n12864 a_23072_n13432.t39 VSS.t499 VSS.t498 nfet_06v0 ad=43.199997f pd=0.6u as=0.2016p ps=1.48u w=0.36u l=0.6u
X1035 a_25544_n16412 a_25573_n12167 VDD.t2100 VDD.t2099 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X1036 a_33440_n2272 a_33292_n2716 a_33272_n2272 VSS.t1517 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
D30 VSS.t680 a_21692_n6694.t10 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1037 VDD.t3227 a_23484_n20052 a_23396_n20008 VDD.t3226 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1038 VDD.t4049 a_44988_n20485 a_44900_n20388 VDD.t4048 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1039 a_13501_n22528.t17 a_11023_n22908.t25 a_11087_n23528.t11 VDD.t208 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1040 VDD.t2128 a_40620_n9509 a_40532_n9412 VDD.t2127 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1041 VDD.t3211 a_43868_n20485 a_43780_n20388 VDD.t3210 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1042 VDD.t3585 a_34012_n16916 a_33924_n16872 VDD.t3584 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1043 VSS.t3735 a_33467_1116 a_30732_332.t0 VSS.t3734 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1044 a_42636_n11077 a_42548_n10980 VSS.t4017 VSS.t4016 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1045 a_30500_n10980 a_23072_n13432.t40 VDD.t493 VDD.t492 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X1046 VDD.t495 a_23072_n13432.t41 a_26635_n12996 VDD.t494 pfet_06v0 ad=0.29465p pd=1.74u as=0.26p ps=1.52u w=1u l=0.5u
X1047 a_34460_n20485 a_34372_n20388 VSS.t2325 VSS.t2324 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1048 a_35244_n15348 a_35156_n15304 VSS.t3144 VSS.t1491 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1049 VDD.t1710 a_42157_n660 a_42277_n1192 VDD.t1709 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1050 VDD.t1051 a_33494_n9860 a_21916_n6694.t1 VDD.t1050 pfet_06v0 ad=0.4941p pd=2.03u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1051 a_25573_n12167 a_24569_n11820 VDD.t3693 VDD.t3692 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1052 a_22588_n16916 a_22500_n16872 VSS.t3450 VSS.t3022 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D31 VSS.t500 a_23072_n13432.t42 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1053 a_37372_n20052 a_37284_n20008 VSS.t2033 VSS.t2032 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1054 VDD.t3726 a_41628_n20485 a_41540_n20388 VDD.t3725 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1055 a_23564_n17700 a_28568_n16066 VDD.t4196 VDD.t4195 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1056 a_33004_n15348 a_32916_n15304 VSS.t1508 VSS.t1507 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1057 a_39357_n2228 a_37221_n3543 VSS.t3546 VSS.t3545 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1058 VDD.t4110 a_25940_n17606.t3 a_26172_n14564.t0 VDD.t4109 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1059 a_36252_n20052 a_36164_n20008 VSS.t2168 VSS.t2167 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1060 a_42972_n1236 a_42884_n1192 VSS.t2253 VSS.t2252 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1061 a_31461_n8248 a_31341_n8292 VSS.t4050 VSS.t4049 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X1062 a_11087_n20850.t27 a_13623_n20230.t22 a_13501_n19850.t17 VSS.t619 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1063 a_31100_n20485 a_31012_n20388 VSS.t3359 VSS.t3358 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1064 a_11087_n23528.t35 a_2167_3472.t67 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X1065 VDD.t2777 a_36140_n15348 a_36052_n15304 VDD.t2776 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1066 VDD.t1264 a_21804_n2273.t3 a_21716_n2229 VDD.t1263 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1067 a_45324_n4805 a_45236_n4708 VSS.t3783 VSS.t3782 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1068 VDD.t2881 a_27597_n8292 a_27717_n7672 VDD.t2880 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1069 VDD.t3313 a_21692_n18484 a_21604_n18440 VDD.t908 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1070 a_25612_n878.t0 a_34953_n1572 VDD.t2820 VDD.t2819 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1071 a_30808_n6334 a_30320_n6636 a_31068_n6276 VDD.t1968 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1072 a_34012_n20052 a_33924_n20008 VSS.t2887 VSS.t2886 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1073 a_43980_n18917 a_43892_n18820 VSS.t4329 VSS.t4328 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1074 a_24913_864 a_22724_860.t2 a_24041_816 VDD.t860 pfet_06v0 ad=0.1079p pd=0.935u as=0.27805p ps=2.17u w=0.415u l=0.5u
X1075 VSS.t936 a_31011_n8292 a_30396_n7508 VSS.t935 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1076 VDD.t3715 a_24088_n16087 a_23564_n20836 VDD.t3714 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1077 VDD.t3174 a_47564_n6373 a_47476_n6276 VDD.t3173 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1078 a_33518_n11592 a_32854_n12168 VSS.t2923 VSS.t2922 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1079 a_41740_n18917 a_41652_n18820 VSS.t2058 VSS.t2057 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1080 a_25936_1564 a_25524_1243 VSS.t1418 VSS.t1417 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1081 a_28352_n320 a_26736_n364 a_27224_n62 VSS.t1527 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1082 VDD.t3207 a_47564_n3237 a_47476_n3140 VDD.t3206 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1083 VDD.t690 a_29800_n5940.t9 a_28156_n6412.t14 VDD.t689 pfet_06v0 ad=0.367p pd=1.92u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1084 a_40620_n18917 a_40532_n18820 VSS.t2060 VSS.t2059 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1085 a_21892_n9816 a_22220_n9860 a_21872_n9394 VSS.t1138 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1086 a_33999_n1400 a_33375_n1976 a_33831_n1400 VDD.t1953 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1087 OUT[0].t3 a_29408_1944.t12 VSS.t3987 VSS.t3986 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1088 VSS.t660 a_21772_1116.t6 a_13623_n4162.t7 VSS.t464 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1089 VDD.t832 a_33776_n5896.t11 a_34708_n5896.t13 VDD.t831 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1090 a_44640_1944.t7 a_44004_n1192 VDD.t2502 VDD.t2501 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1091 VDD.t3225 a_24631_n3588 a_31636_n2760 VDD.t3224 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1092 a_11023_n4162.t18 a_13623_n4162.t20 VDD.t554 VDD.t553 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1093 VDD.t2215 a_46220_n11077 a_46132_n10980 VDD.t2214 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1094 a_25836_n1236.t2 a_34649_n2412 VSS.t3707 VSS.t3706 nfet_06v0 ad=0.2119p pd=1.335u as=0.2119p ps=1.335u w=0.815u l=0.6u
X1095 VSS.t3035 a_33608_n4284 a_33416_n4240 VSS.t3034 nfet_06v0 ad=0.2016p pd=1.48u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1096 a_22364_n10512 a_22264_n10556 VSS.t2263 VSS.t2262 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1097 VDD.t2959 a_44092_n18484 a_44004_n18440 VDD.t2958 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1098 a_28454_n2424 a_28940_n2406.t3 VSS.t3796 VSS.t3795 nfet_06v0 ad=0.3608p pd=2.52u as=0.2911p ps=1.53u w=0.82u l=0.6u
X1099 a_31548_n10172.t14 a_33496_n8222.t11 VDD.t288 VDD.t287 pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1100 a_32732_n10556 a_32424_n10512 VDD.t4180 VDD.t4179 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X1101 a_10778_2852.t0 a_10712_4516.t34 VSS.t339 VSS.t338 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X1102 a_22016_n4257 a_21604_n3844 VDD.t1717 VDD.t1716 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X1103 a_45212_n5940 a_45124_n5896 VSS.t3216 VSS.t3215 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1104 VDD.t4283 a_48012_n9509 a_47924_n9412 VDD.t4282 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1105 a_41392_1944.t5 a_40196_1944 VDD.t3060 VDD.t3059 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1106 VSS.t4199 a_32108_n2332.t18 a_41204_1243 VSS.t4198 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1107 a_35916_n4 a_35816_n174 VSS.t3386 VSS.t3385 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1108 VDD.t2957 a_45772_n101 a_45684_n4 VDD.t2956 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1109 VDD.t3115 a_27055_n1192 a_27511_n1170 VDD.t3114 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1110 a_33496_n6659.t3 CLK.t5 VDD.t1819 VDD.t1818 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X1111 a_11023_n17552.t18 a_13623_n17552.t22 VDD.t90 VDD.t89 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1112 VDD.t1593 a_21772_n452.t7 a_13623_n22908.t3 VDD.t1592 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1113 a_29308_n20485 a_29220_n20388 VSS.t4086 VSS.t4085 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1114 VDD.t1934 a_23036_n16916 a_22948_n16872 VDD.t1933 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1115 VDD.t92 a_13623_n17552.t23 a_11023_n17552.t17 VDD.t91 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1116 a_42636_n9509 a_42548_n9412 VSS.t3090 VSS.t3089 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1117 a_24128_n704 a_22016_n1121 a_23816_n704 VDD.t3362 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X1118 a_24693_n6104 a_24573_n6724 a_23949_n6724 VDD.t2568 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1119 a_44005_n408 a_43885_n452 VSS.t4222 VSS.t4221 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X1120 a_23999_n2320.t1 a_24233_n844 VDD.t3543 VDD.t3542 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1121 a_38716_n4805 a_38628_n4708 VSS.t3366 VSS.t3365 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1122 VDD.t2465 a_27820_n16432 a_27192_n14286 VDD.t2464 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1123 a_26755_n16132 a_27085_n16132 a_27205_n15534 VDD.t1883 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1124 VDD.t4221 a_43555_n452 a_41864_1394 VDD.t4220 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1125 VSS.t2423 a_22444_2253.t10 a_n263_3472.t7 VSS.t2422 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1126 a_25276_n20052 a_25188_n20008 VSS.t4096 VSS.t4095 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1127 VDD.t4281 a_46668_n15781 a_46580_n15684 VDD.t4280 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1128 a_41964_1564 a_41864_1394 VSS.t3962 VSS.t3961 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1129 a_27744_n12908 a_21692_n13308.t18 VSS.t2675 VSS.t2674 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1130 a_23404_816 a_25836_n1236.t10 a_25732_n1192 VDD.t1074 pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1131 VDD.t1746 a_13623_n12196.t24 a_11023_n12196.t5 VDD.t1745 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1132 a_25573_n12167 a_24569_n11820 VSS.t3769 VSS.t3768 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
D32 a_21692_n6694.t11 VDD.t636 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1133 VDD.t2801 a_46668_n12645 a_46580_n12548 VDD.t2800 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1134 a_38828_n18917 a_38740_n18820 VSS.t3445 VSS.t3444 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1135 a_22116_n12548 a_21996_n12996.t5 a_21872_n12530 VDD.t3486 pfet_06v0 ad=0.3172p pd=1.74u as=0.4248p ps=1.94u w=1.22u l=0.5u
X1136 a_37260_n12645 a_37172_n12548 VSS.t3312 VSS.t3311 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1137 a_23036_n20052 a_22948_n20008 VSS.t3013 VSS.t3012 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1138 VDD.t1974 a_23816_n704 a_24233_n844 VDD.t1973 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X1139 VDD.t622 a_28156_n6412.t19 a_26328_n6654.t6 VDD.t621 pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X1140 VDD.t3882 a_44428_n15781 a_44340_n15684 VDD.t3881 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1141 a_26495_n2272 a_23072_n13432.t43 a_25895_n2624 VSS.t501 nfet_06v0 ad=86.399994f pd=0.84u as=0.1989p ps=1.465u w=0.36u l=0.6u
X1142 VDD.t3010 a_40396_n6373 a_40308_n6276 VDD.t3009 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1143 a_31884_n18917 a_31796_n18820 VSS.t3427 VSS.t3426 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1144 VDD.t1621 a_44428_n12645 a_44340_n12548 VDD.t1620 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1145 a_11023_n14874.t4 a_13623_n14874.t23 VDD.t1304 VDD.t1303 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1146 VSS.t2863 a_22588_n2020 a_22500_n1976 VSS.t2862 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1147 VDD.t3317 a_40396_n3237 a_40308_n3140 VDD.t3316 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1148 a_40956_n9076 a_40868_n9032 VSS.t1426 VSS.t1425 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1149 a_35020_n12645 a_34932_n12548 VSS.t2854 VSS.t2853 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1150 a_24481_761.t1 a_30192_n15304.t10 VDD.t2286 VDD.t2285 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1151 VDD.t1306 a_13623_n14874.t24 a_11023_n14874.t5 VDD.t1305 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1152 VDD.t3587 a_37484_n11077 a_37396_n10980 VDD.t3586 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1153 VSS.t1766 a_24752_n16132 a_23564_n8292 VSS.t1765 nfet_06v0 ad=0.2344p pd=1.56u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1154 a_28524_n17349 a_28436_n17252 VSS.t3357 VSS.t2184 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1155 a_26935_n2272 a_25895_n2624 VSS.t3721 VSS.t3720 nfet_06v0 ad=62.1f pd=0.705u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1156 VSS.t558 a_11023_n9518.t24 a_11087_n10138.t4 VSS.t70 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1157 a_41852_n13780 a_41764_n13736 VSS.t3842 VSS.t3841 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1158 a_13623_n17552.t15 a_21772_n8292.t11 VDD.t417 VDD.t416 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1159 VDD.t2830 a_47900_n15348 a_47812_n15304 VDD.t2829 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1160 a_23024_n8544 a_22876_n8988 a_22856_n8544 VSS.t3266 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1161 a_11087_n10138.t5 a_11023_n9518.t25 VSS.t559 VSS.t72 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X1162 a_41852_n10644 a_41764_n10600 VSS.t1282 VSS.t1281 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1163 a_10778_2852.t2 a_10712_4516.t35 VSS.t341 VSS.t340 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1164 a_44629_n408 a_44509_n452 a_43885_n452 VSS.t1317 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X1165 VSS.t127 a_26553_377.t3 a_26431_n1192 VSS.t126 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X1166 VSS.t778 a_24481_761.t29 a_35008_n3456 VSS.t777 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1167 a_33497_n9032 a_32767_n9010 VSS.t1167 VSS.t1166 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X1168 VDD.t3078 a_33686_n11592 a_34142_n12146 VDD.t3077 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1169 a_23024_n5408 a_22876_n5852 a_22856_n5408 VSS.t3079 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1170 a_39612_n12212 a_39524_n12168 VSS.t2784 VSS.t2783 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1171 VDD.t4081 a_35456_n4628.t11 a_32108_n2332.t15 VDD.t4080 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1172 a_45772_n4805 a_45684_n4708 VSS.t2068 VSS.t2067 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1173 a_29940_n8548 a_21916_n6694.t3 a_29736_n8548 VSS.t3900 nfet_06v0 ad=0.1312p pd=1.14u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1174 a_32375_n9032 a_31919_n9032 VDD.t2146 VDD.t2145 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1175 a_23703_n5156.t0 a_28454_n2424 VSS.t3343 VSS.t3342 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1176 a_28764_n8247 a_29123_n6679 a_29176_n7819 VDD.t2532 pfet_06v0 ad=0.4012p pd=1.85u as=0.58035p ps=2.155u w=1.095u l=0.5u
X1177 VDD.t2704 a_38380_n17349 a_38292_n17252 VDD.t2703 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1178 VDD.t3253 a_38380_n14213 a_38292_n14116 VDD.t3252 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1179 a_34649_n2412 a_34232_n2272 a_35025_n2272 VSS.t1023 nfet_06v0 ad=0.3586p pd=2.51u as=0.217p ps=1.515u w=0.815u l=0.6u
X1180 a_38268_n7508 a_38180_n7464 VSS.t1150 VSS.t1149 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1181 a_29900_n10600.t1 a_29444_n10116 VDD.t1964 VDD.t1963 pfet_06v0 ad=0.5368p pd=3.32u as=0.35315p ps=1.96u w=1.22u l=0.5u
X1182 a_45212_332 a_45124_376 VSS.t3188 VSS.t3187 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1183 a_24464_n11680 a_21940_n11684 a_24152_n11680 VSS.t2275 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1184 VDD.t1976 a_36140_n17349 a_36052_n17252 VDD.t1975 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1185 a_23932_n16916 a_23844_n16872 VSS.t2490 VSS.t2489 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1186 a_22876_n4284 a_22568_n4240 VDD.t2971 VDD.t2970 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X1187 VDD.t2876 a_36140_n14213 a_36052_n14116 VDD.t2266 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1188 a_7119_4292 a_1955_4292.t2 VDD.t2352 VDD.t2351 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X1189 a_7119_4292 a_4001_4292.t6 a_3935_4156.t1 VDD.t843 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X1190 a_42948_n1976 a_42244_n1572 VDD.t3798 VDD.t3797 pfet_06v0 ad=0.3477p pd=1.79u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1191 a_31459_n12996 a_31789_n12996 a_31909_n12952 VSS.t4361 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X1192 a_25160_n14816 a_23360_n15233 a_24220_n15260 VSS.t1514 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1193 VSS.t1286 a_37632_n2020 a_25019_n3588.t0 VSS.t1285 nfet_06v0 ad=0.2344p pd=1.56u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1194 a_21692_n6694.t1 a_30900_n9032 VDD.t3678 VDD.t3677 pfet_06v0 ad=0.3782p pd=1.84u as=0.4941p ps=2.03u w=1.22u l=0.5u
X1195 VSS.t780 a_24481_761.t30 a_32880_n10112 VSS.t779 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1196 VDD.t4194 a_28568_n16066 a_23564_n17700 VDD.t4193 pfet_06v0 ad=0.458p pd=2.02u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1197 a_26115_n328 a_25975_n184 a_25627_n452 VSS.t1407 nfet_06v0 ad=0.134p pd=1.1u as=0.176p ps=1.68u w=0.4u l=0.6u
X1198 VDD.t2963 a_47452_n10644 a_47364_n10600 VDD.t2962 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1199 a_45660_n5940 a_45572_n5896 VSS.t3337 VSS.t3336 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1200 a_33292_n2716 a_32984_n2672 VSS.t2049 VSS.t2048 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X1201 VSS.t286 a_31548_n10172.t19 a_33588_n3461 VSS.t285 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1202 VSS.t4349 a_30472_n9815 a_25724_n14564 VSS.t4348 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X1203 a_34895_376 a_34271_376 a_34747_952 VSS.t3532 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1204 VDD.t2549 a_45212_n1669 a_45124_n1572 VDD.t2548 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1205 VDD.t1629 a_45212_n10644 a_45124_n10600 VDD.t1628 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1206 a_25767_n12951 a_24964_n14116 VSS.t1913 VSS.t1912 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1207 a_34908_n18484 a_34820_n18440 VSS.t3252 VSS.t3251 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1208 VDD.t1174 a_23564_n8292 a_21772_n8292.t5 VDD.t1173 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1209 VDD.t3824 a_21916_n6694.t4 a_28736_n4633.t19 VDD.t3823 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X1210 VSS.t3407 a_33488_n12996 a_23564_n14564.t0 VSS.t3406 nfet_06v0 ad=0.2344p pd=1.56u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1211 VSS.t3989 a_29408_1944.t13 OUT[0].t2 VSS.t3988 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1212 a_13623_n4162.t6 a_21772_1116.t7 VSS.t664 VSS.t663 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1213 a_35632_1248 a_24481_761.t31 VSS.t782 VSS.t781 nfet_06v0 ad=43.199997f pd=0.6u as=0.2016p ps=1.48u w=0.36u l=0.6u
X1214 a_34953_n1572 a_34223_n1976 VDD.t2320 VDD.t2319 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X1215 a_32856_n7376 a_32560_n7020 a_31799_n7508 VDD.t1197 pfet_06v0 ad=0.2424p pd=1.465u as=0.25375p ps=1.51u w=0.505u l=0.5u
X1216 VDD.t2869 a_46108_n9076 a_46020_n9032 VDD.t2868 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1217 a_47452_n16916 a_47364_n16872 VSS.t2527 VSS.t2526 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1218 a_47004_n2804 a_46916_n2760 VSS.t4113 VSS.t2231 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1219 VDD.t328 a_10712_4516.t36 a_10778_2852.t3 VDD.t327 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1220 a_30224_376 a_28492_332 VDD.t1363 VDD.t1362 pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1221 a_45212_n16916 a_45124_n16872 VSS.t4276 VSS.t4275 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1222 VDD.t1693 a_37024_1944.t11 OUT[2].t12 VDD.t1692 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1223 VDD.t2287 a_30192_n15304.t11 a_24481_761.t2 VDD.t1648 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1224 VDD.t1379 a_41392_1944.t11 OUT[4].t12 VDD.t1378 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1225 a_32108_n2332.t14 a_35456_n4628.t12 VDD.t4083 VDD.t4082 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1226 a_31628_n5940.t11 a_33496_n6659.t15 VSS.t150 VSS.t149 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X1227 a_44428_n6373 a_44340_n6276 VSS.t3174 VSS.t3173 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1228 a_41740_n3237 a_41652_n3140 VSS.t3165 VSS.t3164 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1229 a_38984_n1975 a_23999_n2320.t2 VSS.t2497 VSS.t2496 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X1230 a_42188_n18917 a_42100_n18820 VSS.t3526 VSS.t3525 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1231 a_37221_n3543 a_36217_n3500 VDD.t1152 VDD.t1151 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1232 VDD.t1792 a_23036_n15781 a_22948_n15684 VDD.t1791 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1233 a_11087_n15494.t27 a_11023_n14874.t24 VSS.t59 VSS.t58 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1234 VDD.t2791 a_39948_n7941 a_39860_n7844 VDD.t2790 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1235 a_22568_n10512 a_21604_n10116 a_22364_n10512 VSS.t3449 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1236 a_22444_332.t0 a_29920_n3900.t11 VDD.t602 VDD.t601 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1237 a_25860_n9032 a_25412_n8501 VDD.t1426 VDD.t1425 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X1238 VSS.t3675 a_27852_n14990 a_27316_n14820 VSS.t3674 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1239 a_31324_n4372 a_31348_n1931 VSS.t1148 VSS.t1147 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X1240 a_29980_n20052 a_29892_n20008 VSS.t2492 VSS.t2491 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1241 a_11023_n20230.t7 a_13623_n20230.t23 VSS.t621 VSS.t620 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1242 a_28860_n20052 a_28772_n20008 VSS.t4129 VSS.t4128 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1243 a_30192_n15304.t1 a_27988_n20388 VSS.t2811 VSS.t2810 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1244 a_36155_n10116 a_30871_n11728 a_33900_n11428 VSS.t958 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1245 VSS.t209 a_13623_n22908.t14 a_11023_n22908.t7 VSS.t208 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X1246 a_26944_n14116 a_26532_n14437 VSS.t2037 VSS.t2036 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1247 VDD.t3886 a_38828_n9509 a_38740_n9412 VDD.t3885 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1248 a_26620_n20052 a_26532_n20008 VSS.t3167 VSS.t3166 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1249 a_11023_n22908.t6 a_13623_n22908.t15 VSS.t211 VSS.t210 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
D33 a_21804_n2273.t4 VDD.t1265 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1250 VSS.t3113 a_29900_760.t6 a_29812_860 VSS.t3112 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1251 VDD.t3752 a_41292_n9509 a_41204_n9412 VDD.t3751 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1252 a_44092_n12212 a_44004_n12168 VSS.t3394 VSS.t3393 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1253 VDD.t3796 a_42244_n1572 a_42948_n1976 VDD.t3795 pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X1254 VSS.t1080 a_30452_n5156.t5 a_27259_804.t0 VSS.t1079 nfet_06v0 ad=0.3608p pd=2.52u as=0.2255p ps=1.37u w=0.82u l=0.6u
X1255 a_30036_n7464 a_29476_n6980 a_29908_n6980 VSS.t2352 nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X1256 VDD.t4085 a_35456_n4628.t13 a_32108_n2332.t13 VDD.t4084 pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1257 VDD.t1034 a_28736_n4633.t20 a_29476_n6980 VDD.t1033 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1258 a_11087_n12816.t7 a_11023_n12196.t24 VSS.t118 VSS.t58 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1259 VDD.t2779 a_37372_n20052 a_37284_n20008 VDD.t2778 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1260 a_32432_n2689 a_32020_n2276 VDD.t3025 VDD.t3024 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X1261 VDD.t2095 a_36252_n20052 a_36164_n20008 VDD.t2094 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1262 a_39276_n9509 a_39188_n9412 VSS.t3350 VSS.t3349 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1263 VDD.t2589 a_24573_n12996 a_24693_n12376 VDD.t2588 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1264 a_11087_n10138.t24 a_13623_n9518.t15 a_13501_n9138.t17 VSS.t245 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1265 a_32628_n10512 a_24481_761.t32 VDD.t724 VDD.t723 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X1266 VDD.t2793 a_34012_n20052 a_33924_n20008 VDD.t2792 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1267 a_35356_n16916 a_35268_n16872 VSS.t1459 VSS.t1458 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1268 VSS.t727 a_13623_n6840.t23 a_11023_n6840.t4 VSS.t726 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1269 a_37499_860 a_25612_n878.t3 a_30104_n1148 VSS.t845 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1270 VDD.t1254 a_31544_1248 a_31961_1204 VDD.t1253 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X1271 a_30451_n452 a_30781_n452 a_30901_146 VDD.t3324 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1272 a_36593_n3456 a_24481_761.t33 VSS.t784 VSS.t783 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X1273 a_33116_n16916 a_33028_n16872 VSS.t1243 VSS.t1242 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1274 a_13501_n6460.t10 a_11023_n6840.t25 a_11087_n7460.t25 VDD.t111 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1275 VDD.t1899 a_34460_n18484 a_34372_n18440 VDD.t1898 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1276 a_44005_146 a_43885_n452 VDD.t4149 VDD.t4148 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X1277 a_25577_n14956 a_25160_n14816 a_25953_n14816 VSS.t1982 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X1278 VDD.t2022 a_137_4292 a_3025_2852 VDD.t2021 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X1279 a_22588_n2020 a_22918_n2020 a_23038_n1976 VSS.t4112 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X1280 VDD.t4249 a_23564_n17700 a_21772_n17700.t7 VDD.t4248 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1281 VDD.t2204 a_32220_n18484 a_32132_n18440 VDD.t2203 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1282 VDD.t3738 a_23564_n14564.t3 a_21772_n14564.t1 VDD.t3737 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1283 a_33653_952 a_33533_908 a_32909_841 VSS.t3127 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X1284 VDD.t3038 a_45660_n1669 a_45572_n1572 VDD.t3037 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1285 a_33496_n8222.t5 a_34708_n5896.t17 VDD.t446 VDD.t445 pfet_06v0 ad=0.2952p pd=1.54u as=0.367p ps=1.92u w=0.82u l=0.5u
X1286 a_37024_1944.t5 a_36388_1944 VDD.t1655 VDD.t1654 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1287 a_13623_n22908.t2 a_21772_n452.t8 VDD.t1595 VDD.t1594 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1288 a_44316_n1236 a_44228_n1192 VSS.t2009 VSS.t2008 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1289 VSS.t3848 a_21692_2431 a_28671_n1976 VSS.t3847 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X1290 a_48012_n4805 a_47924_n4708 VSS.t1892 VSS.t1891 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1291 VDD.t604 a_29920_n3900.t12 a_22444_332.t1 VDD.t603 pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1292 VSS.t860 a_34708_n5896.t18 a_35456_n4628.t2 VSS.t859 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1293 VDD.t3249 a_46556_n9076 a_46468_n9032 VDD.t3248 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1294 a_47452_n2804 a_47364_n2760 VSS.t3666 VSS.t1141 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1295 VSS.t2792 a_22052_1944 a_29408_1944.t1 VSS.t2791 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1296 VDD.t3103 a_46108_n15348 a_46020_n15304 VDD.t3102 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1297 a_10712_4516.t29 a_10778_2852.t18 VDD.t367 VDD.t366 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1298 VSS.t49 a_21772_n8292.t12 a_13623_n17552.t4 VSS.t48 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1299 a_13501_n14494.t17 a_11023_n14874.t25 a_11087_n15494.t17 VDD.t75 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1300 a_22096_376 a_21996_332.t2 VDD.t438 VDD.t437 pfet_06v0 ad=0.4248p pd=1.94u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1301 VDD.t2992 a_39164_n16916 a_39076_n16872 VDD.t2991 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1302 a_11087_n15494.t16 a_11023_n14874.t26 a_13501_n14494.t16 VDD.t76 pfet_03v3 ad=0.728p pd=3.32u as=1.82p ps=6.9u w=2.8u l=0.28u
X1303 a_30104_n1148 a_25612_n878.t4 VDD.t795 VDD.t794 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1304 a_44876_n6373 a_44788_n6276 VSS.t3081 VSS.t3080 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1305 a_39612_n9076 a_39524_n9032 VSS.t3881 VSS.t3880 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1306 VDD.t3930 a_39164_n13780 a_39076_n13736 VDD.t3929 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D34 a_24481_761.t34 VDD.t725 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1307 a_28863_n10116 a_28437_n13705 a_28435_n10599 VSS.t2624 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X1308 a_46668_n11077 a_46580_n10980 VSS.t3507 VSS.t3506 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1309 VDD.t1778 a_35916_n12645 a_35828_n12548 VDD.t1777 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1310 a_25237_n10599 a_24233_n10252 VDD.t993 VDD.t992 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1311 VDD.t2197 a_25276_n20052 a_25188_n20008 VDD.t2196 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1312 a_37372_n20485 a_37284_n20388 VSS.t2913 VSS.t2912 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1313 a_13501_n17172.t16 a_11023_n17552.t26 a_11087_n18172.t16 VDD.t403 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1314 VSS.t786 a_24481_761.t35 a_33440_n2272 VSS.t785 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1315 a_44428_n11077 a_44340_n10980 VSS.t3015 VSS.t3014 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1316 a_36252_n20485 a_36164_n20388 VSS.t3115 VSS.t3114 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1317 a_25137_864 a_22724_860.t3 a_24913_864 VSS.t915 nfet_06v0 ad=0.2898p pd=2.33u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1318 a_46668_n101 a_46580_n4 VSS.t4056 VSS.t4055 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1319 a_34176_n6976 a_32455_n7420 a_33048_n7420 VDD.t4261 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1320 VDD.t2939 a_23036_n20052 a_22948_n20008 VDD.t2938 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1321 EOC.t10 a_45648_1564.t16 VDD.t56 VDD.t55 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1322 a_36576_n320 a_36428_n53 a_36408_n320 VSS.t2859 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1323 a_23619_n12996 a_23949_n12996 a_24069_n12398 VDD.t1192 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1324 a_39164_n20052 a_39076_n20008 VSS.t2111 VSS.t2110 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1325 a_34012_n20485 a_33924_n20388 VSS.t2920 VSS.t2919 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1326 VDD.t2990 a_28232_n12606 a_28040_n12493 VDD.t2989 pfet_06v0 ad=0.2222p pd=1.89u as=0.2424p ps=1.465u w=0.505u l=0.5u
X1327 VSS.t1176 a_25084_1564 a_33216_1944.t3 VSS.t1175 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1328 a_2167_3472.t31 a_11023_n4162.t23 VSS.t2753 VDD.t2691 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1329 a_26531_n8639 a_26861_n8567 a_26981_n9010 VDD.t2926 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1330 a_45324_n9509 a_45236_n9412 VSS.t2858 VSS.t2857 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1331 a_13501_n11816.t7 a_11023_n12196.t25 a_11087_n12816.t17 VDD.t129 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1332 VDD.t3336 a_23484_n18484 a_23396_n18440 VDD.t3335 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1333 a_11087_n12816.t16 a_11023_n12196.t26 a_13501_n11816.t6 VDD.t130 pfet_03v3 ad=0.728p pd=3.32u as=1.82p ps=6.9u w=2.8u l=0.28u
X1334 a_45772_n18917 a_45684_n18820 VSS.t2885 VSS.t2884 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1335 a_11087_n23528.t36 a_2167_3472.t66 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X1336 VSS.t130 a_31628_n5940.t33 a_29800_n5940.t2 VSS.t23 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1337 a_13501_n6460.t3 a_13623_n6840.t24 a_11087_n7460.t3 VSS.t728 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X1338 a_11087_n23528.t37 a_2167_3472.t65 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X1339 a_27134_n13160 a_26470_n13736 VSS.t1268 VSS.t1267 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1340 a_22464_n7393 a_22052_n6980 VSS.t1556 VSS.t1555 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1341 a_43532_n18917 a_43444_n18820 VSS.t3356 VSS.t3355 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1342 a_11087_n18172.t7 a_13623_n17552.t24 a_13501_n17172.t7 VSS.t82 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1343 a_31909_n13966 a_31789_n14564 VDD.t2479 VDD.t2478 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X1344 a_13623_n20230.t5 a_21772_n3588.t8 VSS.t612 VSS.t611 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1345 VDD.t3135 a_43084_n6373 a_42996_n6276 VDD.t3134 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1346 a_29532_n4372.t1 a_21916_n6694.t5 VDD.t3826 VDD.t3825 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1347 a_28644_n9815 a_24348_n16087.t4 VSS.t2513 VSS.t2512 nfet_06v0 ad=0.2119p pd=1.335u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1348 VDD.t1888 a_43084_n3237 a_42996_n3140 VDD.t1887 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1349 VDD.t25 a_24815_n3588.t7 a_28736_n4633.t3 VDD.t24 pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
X1350 a_26702_n9240 a_26266_n9240 a_26470_n9322 VDD.t996 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1351 a_32650_n12168 a_32026_n12168 a_32502_n11592 VSS.t3779 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1352 a_26983_n12728 a_27639_n12537 a_27535_n12493 VDD.t2082 pfet_06v0 ad=0.25375p pd=1.51u as=0.1313p ps=1.025u w=0.505u l=0.5u
X1353 a_10712_4516.t28 a_10778_2852.t19 VDD.t369 VDD.t368 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1354 a_43644_n9076 a_43556_n9032 VSS.t4258 VSS.t4257 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1355 VDD.t2799 a_48012_n11077 a_47924_n10980 VDD.t2798 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1356 a_24385_864 a_23728_464 VSS.t1972 VSS.t1971 nfet_06v0 ad=86.399994f pd=0.84u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1357 VDD.t606 a_29920_n3900.t13 a_33375_n1976 VDD.t605 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1358 a_28048_1248 a_25524_1243 a_27736_1248 VSS.t1416 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1359 a_31292_n2804 a_31324_n4372 VDD.t4027 VDD.t4026 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
D35 a_24481_761.t36 VDD.t726 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1360 a_26859_n3544 a_26383_n2968 a_26607_n3544 VSS.t1702 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X1361 a_23524_464 a_23404_816 VSS.t1637 VSS.t1636 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1362 VDD.t576 a_21772_n3588.t9 a_13623_n20230.t13 VDD.t575 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1363 a_28852_n8292.t0 a_29900_n10600.t3 VDD.t3859 VDD.t3858 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1364 VDD.t2808 a_37820_n10644 a_37732_n10600 VDD.t2807 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1365 a_21692_n15781 a_21604_n15684 VSS.t2926 VSS.t1745 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1366 a_24128_n8544 a_22016_n8961 a_23816_n8544 VDD.t1022 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X1367 VDD.t4069 a_41404_n9076 a_41316_n9032 VDD.t4068 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1368 a_26396_n20485 a_26308_n20388 VSS.t3021 VSS.t3020 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1369 VSS.t2754 a_11023_n4162.t24 VSS.t2754 VSS.t70 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.28u
X1370 a_24128_n5408 a_22016_n5825 a_23816_n5408 VDD.t3073 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
D36 a_25940_n17606.t4 VDD.t4111 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1371 VDD.t1156 a_27190_n5112 a_27646_n4558 VDD.t1155 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1372 a_25237_n5895 a_24233_n5548 VDD.t2953 VDD.t2952 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1373 a_33496_n8222.t4 a_34708_n5896.t19 VDD.t816 VDD.t815 pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X1374 a_42624_1248 a_42476_1515 a_42456_1248 VSS.t4097 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1375 VDD.t670 a_13623_n6840.t25 a_11023_n6840.t5 VDD.t669 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1376 a_24965_n9860 a_21996_n12996.t6 a_25844_n14116 VDD.t3487 pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
D37 a_22140_n6694.t7 VDD.t4060 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1377 VDD.t3545 a_45324_n101 a_45236_n4 VDD.t3544 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1378 a_23319_n2759 a_23999_n2320.t3 VDD.t2407 VDD.t2406 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1379 a_27068_n20052 a_26980_n20008 VSS.t3230 VSS.t3229 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1380 a_37820_n16916 a_37732_n16872 VSS.t2786 VSS.t2785 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1381 a_n263_3472.t13 a_22444_2253.t11 VDD.t2338 VDD.t455 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1382 VSS.t574 a_13623_n4162.t21 a_11023_n4162.t7 VSS.t573 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X1383 a_29532_n4372.t2 a_29900_n10600.t4 VDD.t3861 VDD.t3860 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1384 a_31215_n11684 a_28940_n2406.t4 a_30787_n12167 VSS.t3797 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X1385 a_36700_n16916 a_36612_n16872 VSS.t2595 VSS.t2594 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1386 VDD.t3040 a_23816_n5408 a_24233_n5548 VDD.t3039 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X1387 a_23072_n13432.t1 a_29744_n15604.t13 VSS.t1728 VSS.t1727 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1388 a_23912_n15216 a_23360_n15233 a_23708_n15216 VDD.t1453 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
D38 a_23072_n13432.t44 VDD.t496 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1389 a_29147_n1976 a_28671_n1976 VSS.t3863 VSS.t3862 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1390 a_39052_n12645 a_38964_n12548 VSS.t3178 VSS.t3177 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1391 a_34796_n18917 a_34708_n18820 VSS.t4125 VSS.t4124 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1392 VSS.t1040 a_25237_n10599 a_25642_n9816 VSS.t1039 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X1393 a_41336_n407 a_25539_n407.t2 VDD.t1704 VDD.t1703 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X1394 a_31544_n6592 a_30616_n6221 a_31376_n6592 VSS.t2199 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1395 VDD.t1695 a_37024_1944.t12 OUT[2].t11 VDD.t1694 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1396 VDD.t2202 a_40396_n12645 a_40308_n12548 VDD.t2201 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1397 VSS.t3991 a_29408_1944.t14 OUT[0].t1 VSS.t3990 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1398 a_31436_n18917 a_31348_n18820 VSS.t3232 VSS.t3231 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1399 a_24348_n16087.t0 a_25577_n14956 VSS.t2889 VSS.t2888 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1400 VSS.t3315 a_36520_n3868 a_26388_n17606.t0 VSS.t3314 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X1401 VDD.t3095 a_36773_n5468 a_29612_n8292 VDD.t3094 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1402 VDD.t4200 a_39276_n11077 a_39188_n10980 VDD.t4199 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1403 a_11087_n23528.t38 a_2167_3472.t64 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X1404 a_41852_n18484 a_41764_n18440 VSS.t2323 VSS.t2322 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1405 a_26971_n14820 a_23479_n5156 a_21772_n9860 VSS.t2315 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1406 a_11023_n6840.t6 a_13623_n6840.t26 VSS.t730 VSS.t729 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1407 a_41852_n15348 a_41764_n15304 VSS.t1882 VSS.t1881 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1408 a_43644_n13780 a_43556_n13736 VSS.t2201 VSS.t2200 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1409 a_39948_n3237 a_39860_n3140 VSS.t4131 VSS.t4130 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1410 VSS.t576 a_13623_n4162.t22 a_2167_3472.t1 VSS.t575 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X1411 a_30378_n5112 a_24815_n3588.t8 a_30174_n5112 VSS.t18 nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1412 VDD.t2591 a_37820_n9076 a_37732_n9032 VDD.t2590 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1413 VDD.t3205 a_37036_n11077 a_36948_n10980 VDD.t3204 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1414 VSS.t343 a_10712_4516.t37 a_10778_2852.t4 VSS.t342 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1415 VSS.t3902 a_21916_n6694.t6 a_35595_n8548 VSS.t3901 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1416 a_43644_n10644 a_43556_n10600 VSS.t2331 VSS.t2330 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1417 a_27485_n8500 a_21872_n9394 VDD.t2111 VDD.t955 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1418 a_30092_n10980 a_29992_n11150 VDD.t2949 VDD.t2948 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X1419 VDD.t3356 a_31459_n12996 a_31279_n11728 VDD.t3355 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1420 VDD.t1381 a_41392_1944.t12 OUT[4].t11 VDD.t1380 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1421 a_45772_n9509 a_45684_n9412 VSS.t3228 VSS.t3227 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1422 a_32337_n11296 a_23072_n13432.t45 VSS.t503 VSS.t502 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X1423 a_41404_n13780 a_41316_n13736 VSS.t2632 VSS.t2631 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1424 VDD.t4254 a_29980_n20052 a_29892_n20008 VDD.t4253 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1425 a_41404_n10644 a_41316_n10600 VSS.t3364 VSS.t3363 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1426 a_10712_4516.t16 a_10778_2852.t20 VSS.t379 VSS.t378 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X1427 VDD.t62 a_21692_n5111.t3 a_24628_n363 VDD.t61 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
D39 VSS.t504 a_23072_n13432.t46 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1428 VDD.t4056 a_28860_n20052 a_28772_n20008 VDD.t4055 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1429 VDD.t3506 a_27224_n62 a_27032_51 VDD.t3505 pfet_06v0 ad=0.2222p pd=1.89u as=0.2424p ps=1.465u w=0.505u l=0.5u
X1430 VDD.t3328 a_27452_n2716 a_27348_n2672 VDD.t3327 pfet_06v0 ad=0.22725p pd=1.91u as=0.1313p ps=1.025u w=0.505u l=0.5u
X1431 a_28736_n4633.t2 a_24815_n3588.t9 VDD.t27 VDD.t26 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X1432 a_11087_n18172.t31 a_2167_3472.t79 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X1433 a_41292_n4805 a_41204_n4708 VSS.t3263 VSS.t3262 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1434 a_27535_n12493 a_26635_n12996 VDD.t2060 VDD.t2059 pfet_06v0 ad=0.1313p pd=1.025u as=0.29465p ps=1.74u w=0.505u l=0.5u
X1435 a_24380_n18917 a_24292_n18820 VSS.t3290 VSS.t3289 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1436 a_n263_3472.t6 a_22444_2253.t12 VSS.t2425 VSS.t2424 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1437 VDD.t58 a_45648_1564.t17 EOC.t9 VDD.t57 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1438 a_32984_n2672 a_32020_n2276 a_32780_n2672 VSS.t3109 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1439 a_27001_n4328.t0 a_26271_n4306 VSS.t2915 VSS.t2914 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X1440 a_35456_n4628.t6 a_34708_n5896.t20 VDD.t818 VDD.t817 pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X1441 a_47116_n6373 a_47028_n6276 VSS.t4339 VSS.t4338 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1442 VDD.t3165 a_38380_n18917 a_38292_n18820 VDD.t3164 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1443 a_27485_n8500 a_21872_n9394 VSS.t2190 VSS.t2189 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1444 VDD.t2771 a_26620_n20052 a_26532_n20008 VDD.t2770 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1445 a_21772_n3588.t0 a_23564_n3588.t2 VSS.t2989 VSS.t2988 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1446 a_23816_n3840 a_22016_n4257 a_22876_n4284 VSS.t3352 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1447 a_22140_n18917 a_22052_n18820 VSS.t2194 VSS.t2193 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1448 VDD.t3306 a_36140_n18917 a_36052_n18820 VDD.t3305 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1449 a_32780_n2672 a_31392_n2760 VDD.t4146 VDD.t4145 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X1450 a_29744_n15604.t1 a_24481_761.t37 VSS.t788 VSS.t787 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1451 a_29800_n5940.t1 a_31628_n5940.t34 VSS.t132 VSS.t131 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1452 a_30296_n10980 a_29744_n10980 a_30092_n10980 VDD.t3583 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1453 a_37844_1564 a_37396_1205 VDD.t2769 VDD.t2768 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X1454 a_43845_376 a_43725_908 a_43101_841 VDD.t2108 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1455 a_26006_n5112 a_25530_n5112 VSS.t3840 VSS.t3839 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1456 VSS.t2015 a_37859_377 a_39868_n408 VSS.t2014 nfet_06v0 ad=0.2132p pd=1.34u as=98.399994f ps=1.06u w=0.82u l=0.6u
X1457 VSS.t2677 a_21692_n13308.t19 a_21604_n8548 VSS.t2676 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1458 VSS.t1036 a_24233_n10252 a_24128_n10112 VSS.t1035 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X1459 a_22564_n5112 a_22444_n5156 VSS.t2591 VSS.t2590 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1460 a_21692_n13308.t4 a_26328_n6654.t14 VSS.t2667 VSS.t2666 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1461 VDD.t2871 a_47004_n10644 a_46916_n10600 VDD.t2870 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1462 a_25844_n14116 a_25724_n14564 VDD.t2969 VDD.t2968 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X1463 VDD.t3434 a_28153_1204 a_28048_1248 VDD.t3433 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X1464 a_34272_n4 a_33508_n408 a_34068_n4 VDD.t4262 pfet_06v0 ad=0.4758p pd=2u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1465 a_27628_n3841 a_24815_n3588.t10 VSS.t20 VSS.t19 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X1466 VDD.t3143 a_41852_n9076 a_41764_n9032 VDD.t3142 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1467 a_30876_n18484 a_30788_n18440 VSS.t2962 VSS.t2961 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1468 a_47004_n7508 a_46916_n7464 VSS.t2105 VSS.t2104 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1469 VDD.t3575 a_40060_n10644 a_39972_n10600 VDD.t3574 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1470 VSS.t345 a_10712_4516.t38 a_10778_2852.t5 VSS.t344 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
D40 VSS.t681 a_21692_n6694.t12 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1471 a_24752_n8292 a_25020_n8200.t2 VSS.t900 VSS.t899 nfet_06v0 ad=0.1584p pd=1.6u as=0.2344p ps=1.56u w=0.36u l=0.6u
X1472 VDD.t2403 a_38716_n15348 a_38628_n15304 VDD.t2402 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1473 a_31405_n452 a_22672_n2214.t3 VDD.t1447 VDD.t1446 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1474 a_28247_n10599 a_28519_n10160.t5 a_28435_n10599 VDD.t787 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1475 VSS.t560 a_11023_n9518.t26 a_11087_n10138.t6 VSS.t54 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1476 VSS.t288 a_31548_n10172.t20 a_31460_n10116 VSS.t287 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1477 a_47004_n16916 a_46916_n16872 VSS.t2183 VSS.t2182 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1478 a_28156_n6412.t13 a_29800_n5940.t10 VDD.t696 VDD.t695 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1479 VSS.t1354 a_13623_n14874.t25 a_11023_n14874.t6 VSS.t1353 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1480 a_23708_n15216 a_23608_n15260 VSS.t3388 VSS.t3387 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1481 VDD.t371 a_10778_2852.t21 a_10712_4516.t27 VDD.t370 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1482 VSS.t22 a_24815_n3588.t11 a_34736_n3840 VSS.t21 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1483 VDD.t3020 a_32073_n844 a_31968_n704 VDD.t3019 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X1484 a_33120_n3884 a_32108_n2332.t19 VDD.t4128 VDD.t4127 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X1485 a_40060_n16916 a_39972_n16872 VSS.t2043 VSS.t2042 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1486 a_28352_n320 a_26631_7 a_27224_n62 VDD.t1430 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1487 VDD.t29 a_24815_n3588.t12 a_24731_n3124.t0 VDD.t28 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1488 a_28568_n16066 a_28752_n15348 VDD.t3126 VDD.t3125 pfet_06v0 ad=0.4488p pd=2.92u as=0.458p ps=2.02u w=1.02u l=0.5u
X1489 VSS.t666 a_28156_n6412.t20 a_26440_n5940.t2 VSS.t665 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1490 a_33494_n9860 a_28519_n10160.t6 VSS.t843 VSS.t842 nfet_06v0 ad=0.3608p pd=2.52u as=0.2911p ps=1.53u w=0.82u l=0.6u
X1491 a_28040_n12493 a_27744_n12908 a_26983_n12728 VDD.t1504 pfet_06v0 ad=0.2424p pd=1.465u as=0.25375p ps=1.51u w=0.505u l=0.5u
X1492 a_10778_2852.t10 a_4001_4292.t7 VSS.t890 VSS.t348 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1493 a_28524_n18484 a_28436_n18440 VSS.t2185 VSS.t2184 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1494 a_25544_n16412 a_25573_n12167 VSS.t2170 VSS.t2169 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X1495 VDD.t3342 a_46668_n7941 a_46580_n7844 VDD.t3341 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1496 VDD.t3201 a_28076_n17349 a_27988_n17252 VDD.t3200 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1497 VDD.t2135 a_46668_n4805 a_46580_n4708 VDD.t2134 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1498 a_40620_n9509 a_40532_n9412 VSS.t2205 VSS.t2204 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1499 a_26563_n12212 a_27404_n14990 a_27316_n14820 VSS.t3360 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1500 VDD.t2339 a_22444_2253.t13 a_n263_3472.t12 VDD.t459 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1501 VDD.t3130 a_39164_n7508 a_39076_n7464 VDD.t3129 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1502 VDD.t2087 a_34908_n20485 a_34820_n20388 VDD.t2086 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1503 a_34403_332 a_34068_n4 VSS.t1933 VSS.t1932 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1504 a_44509_n452 a_42948_n1976 VSS.t3070 VSS.t3069 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1505 a_25500_n20485 a_25412_n20388 VSS.t3205 VSS.t3204 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1506 VSS.t2790 a_22052_1944 a_29408_1944.t0 VSS.t2789 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1507 VDD.t2802 a_39164_n4372 a_39076_n4328 VDD.t2794 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1508 a_29532_n20052 a_29444_n20008 VSS.t3973 VSS.t3972 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1509 a_22772_n13648 a_23072_n13432.t47 VDD.t498 VDD.t497 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X1510 a_27337_n3140 a_26607_n3544 VSS.t4300 VSS.t4299 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X1511 a_45324_n101 a_45236_n4 VSS.t4347 VSS.t4346 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1512 a_29800_n5940.t5 a_31628_n5940.t35 VDD.t142 VDD.t141 pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X1513 VDD.t3987 a_38268_n10644 a_38180_n10600 VDD.t3986 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1514 VSS.t1830 a_13623_n12196.t25 a_11023_n12196.t6 VSS.t1829 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1515 a_28412_n20052 a_28324_n20008 VSS.t1993 VSS.t1992 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1516 a_30372_376 a_29900_760.t7 a_30224_376 VDD.t2222 pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X1517 a_11023_n17552.t6 a_13623_n17552.t25 VSS.t84 VSS.t83 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1518 VSS.t4181 a_25940_n17606.t5 a_25600_n5895 VSS.t4180 nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
X1519 a_24573_n6724 a_22544_n4690 VSS.t2091 VSS.t2090 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1520 VDD.t2840 a_43980_n15781 a_43892_n15684 VDD.t2839 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1521 VSS.t3491 a_23564_1116.t3 a_21772_1116.t1 VSS.t3490 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1522 a_27485_n10068 a_25573_n12167 VDD.t2098 VDD.t2097 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1523 VDD.t3870 a_39164_n20052 a_39076_n20008 VDD.t986 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D41 a_26388_n17606.t4 VDD.t205 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1524 a_24233_n844 a_23816_n704 a_24609_n704 VSS.t2050 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X1525 a_30296_n10980 a_29332_n11301 a_30092_n10980 VSS.t3557 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1526 VDD.t3948 a_43980_n12645 a_43892_n12548 VDD.t3947 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1527 VDD.t3006 a_41740_n15781 a_41652_n15684 VDD.t3005 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1528 a_34727_376 a_34271_376 VDD.t3448 VDD.t3447 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1529 VDD.t728 a_24481_761.t38 a_31451_n7508 VDD.t727 pfet_06v0 ad=0.29465p pd=1.74u as=0.26p ps=1.52u w=1u l=0.5u
X1530 a_24041_816 a_23728_464 VDD.t1897 VDD.t1896 pfet_06v0 ad=0.1521p pd=1.105u as=0.3975p ps=2.185u w=0.585u l=0.5u
X1531 a_24681_n7116 a_23072_n13432.t48 VDD.t500 VDD.t499 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X1532 VDD.t3163 a_41740_n12645 a_41652_n12548 VDD.t3162 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1533 a_33900_n18917 a_33812_n18820 VSS.t3855 VSS.t3854 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1534 a_38268_n16916 a_38180_n16872 VSS.t1808 VSS.t1807 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1535 VDD.t3153 a_40620_n15781 a_40532_n15684 VDD.t3152 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1536 a_26383_n2968 a_25759_n3544 a_26235_n3544 VSS.t3570 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1537 a_47564_n6373 a_47476_n6276 VSS.t2893 VSS.t2892 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1538 OUT[4].t10 a_41392_1944.t13 VDD.t1383 VDD.t1382 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1539 a_35816_n174 a_35119_398 VSS.t435 VSS.t434 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X1540 a_23192_n11680 a_22352_n12097 a_22904_n12080 VSS.t1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1541 a_26235_2520 a_25759_1944 VSS.t951 VSS.t950 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1542 VSS.t3600 a_30584_n1954 a_21996_n12996.t1 VSS.t3599 nfet_06v0 ad=0.151p pd=1.185u as=0.1261p ps=1.005u w=0.485u l=0.6u
X1543 VDD.t3936 a_37372_n18484 a_37284_n18440 VDD.t3935 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1544 a_44876_n15781 a_44788_n15684 VSS.t3960 VSS.t3959 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1545 a_11023_n20230.t6 a_13623_n20230.t24 VSS.t623 VSS.t622 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1546 VDD.t3828 a_36252_n18484 a_36164_n18440 VDD.t3827 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1547 VDD.t3467 a_33672_n10112 a_34089_n10252 VDD.t3466 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X1548 VSS.t2179 a_34895_376 a_35371_951 VSS.t2178 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X1549 VDD.t608 a_29920_n3900.t14 a_24815_n3588.t3 VDD.t607 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1550 VSS.t1817 a_27485_n10068 a_27605_n10024 VSS.t1816 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1551 a_42636_n15781 a_42548_n15684 VSS.t1771 VSS.t1770 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1552 a_22564_n5112 a_22892_n5156.t3 a_22544_n4690 VSS.t4215 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1553 a_48012_n9509 a_47924_n9412 VSS.t3398 VSS.t3397 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1554 VDD.t1281 a_34012_n18484 a_33924_n18440 VDD.t1280 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1555 a_21692_n13308.t3 a_26328_n6654.t15 VSS.t2669 VSS.t2668 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1556 VDD.t1340 a_43196_n7508 a_43108_n7464 VDD.t1339 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1557 VDD.t3914 a_43196_n4372 a_43108_n4328 VDD.t3913 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1558 a_28435_n10599 a_28335_n10644 a_28247_n10599 VDD.t1092 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1559 a_30575_n2276 a_22220_690.t7 VSS.t834 VSS.t833 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1560 a_47452_n7508 a_47364_n7464 VSS.t2985 VSS.t2984 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1561 a_37585_n3140 a_22052_n4708 VDD.t3609 VDD.t3608 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1562 VDD.t3550 a_43308_n5940 a_43220_n5896 VDD.t3549 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1563 a_21916_n6694.t0 a_33494_n9860 VSS.t1088 VSS.t1087 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1564 a_29540_n11728 a_26388_n17606.t5 VSS.t233 VSS.t232 nfet_06v0 ad=0.14p pd=1.1u as=0.224p ps=1.52u w=0.4u l=0.6u
X1565 VDD.t3843 a_43196_n15348 a_43108_n15304 VDD.t3842 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1566 VDD.t3833 a_39948_n12645 a_39860_n12548 VDD.t3832 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1567 VDD.t972 a_38828_n15781 a_38740_n15684 VDD.t971 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1568 a_33940_n408 a_33820_n452.t2 VSS.t3883 VSS.t3882 nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1569 a_28156_n6412.t12 a_29800_n5940.t11 VDD.t698 VDD.t697 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1570 a_11087_n23528.t39 a_2167_3472.t63 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X1571 a_33029_398 a_32909_841 VDD.t4252 VDD.t4251 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X1572 a_34747_n616 a_34271_n1192 VSS.t1404 VSS.t1403 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1573 VDD.t1723 a_45212_n7508 a_45124_n7464 VDD.t1722 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1574 VDD.t985 a_37708_n12645 a_37620_n12548 VDD.t984 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1575 VDD.t3149 a_27068_n20052 a_26980_n20008 VDD.t3148 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1576 VDD.t3847 a_45212_n4372 a_45124_n4328 VDD.t3846 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1577 a_27022_n5112 a_26358_n4618 VSS.t1453 VSS.t1452 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1578 a_30604_n11029 a_30296_n10980 VSS.t4107 VSS.t4106 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
D42 VSS.t1306 a_21804_n2273.t5 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1579 a_40396_n6373 a_40308_n6276 VSS.t2848 VSS.t2847 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1580 a_39164_n20485 a_39076_n20388 VSS.t3911 VSS.t3910 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1581 VSS.t397 a_21692_n5468.t19 a_25524_1243 VSS.t396 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1582 a_40620_n5940 a_40532_n5896 VSS.t2251 VSS.t2250 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1583 a_22364_n4240 a_21792_n7464 VSS.t1067 VSS.t1066 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1584 VSS.t697 a_21772_n20836.t12 a_13623_n6840.t5 VSS.t696 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1585 a_22340_376 a_22220_690.t8 a_22096_376 VDD.t779 pfet_06v0 ad=0.3172p pd=1.74u as=0.4248p ps=1.94u w=1.22u l=0.5u
X1586 a_29744_n10980 a_29332_n11301 VDD.t3476 VDD.t3475 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X1587 a_13623_n6840.t4 a_21772_n20836.t13 VSS.t699 VSS.t698 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1588 a_27709_n16132 a_24348_n16087.t5 VDD.t2429 VDD.t2428 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1589 a_13623_n4162.t5 a_21772_1116.t8 VSS.t556 VSS.t555 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1590 a_39544_420 a_38951_420 a_40280_864 VSS.t3299 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1591 a_11087_n20850.t32 a_2167_3472.t19 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X1592 VDD.t2500 a_44004_n1192 a_44640_1944.t6 VDD.t2499 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1593 VDD.t1936 a_23816_n10112 a_24233_n10252 VDD.t1935 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X1594 a_13501_n19850.t16 a_13623_n20230.t25 a_11087_n20850.t26 VSS.t624 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1595 VDD.t3539 a_25276_n18484 a_25188_n18440 VDD.t3538 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1596 a_34465_n10112 a_24481_761.t39 VSS.t790 VSS.t789 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X1597 VSS.t2844 a_43644_n705 a_43556_n661 VSS.t2843 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1598 a_30616_n3544 a_27259_804.t8 a_22444_332.t4 VSS.t854 nfet_06v0 ad=0.1722p pd=1.24u as=0.4161p ps=1.905u w=0.82u l=0.6u
X1599 VDD.t1697 a_37024_1944.t13 OUT[2].t10 VDD.t1696 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1600 VDD.t1530 a_31787_n3969 a_29920_n3900.t1 VDD.t1529 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1601 a_26154_n4536 a_25530_n5112 a_26006_n5112 VSS.t3838 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1602 VSS.t152 a_33496_n6659.t16 a_31628_n5940.t10 VSS.t151 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X1603 a_11087_n23528.t7 a_13623_n22908.t16 a_13501_n22528.t7 VSS.t212 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1604 a_47564_n18917 a_47476_n18820 VSS.t3905 VSS.t3904 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1605 VDD.t3562 a_23036_n18484 a_22948_n18440 VDD.t3343 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1606 a_25160_n14816 a_22948_n14820 a_24220_n15260 VDD.t937 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X1607 a_37024_1944.t3 a_36388_1944 VSS.t1742 VSS.t1741 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1608 a_29744_n15604.t0 a_24481_761.t40 VSS.t791 VSS.t695 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1609 VSS.t2755 a_11023_n4162.t25 VSS.t2755 VSS.t60 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.28u
X1610 a_45324_n18917 a_45236_n18820 VSS.t4002 VSS.t4001 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1611 a_26742_n13160 a_26266_n13736 a_26470_n13736 VSS.t4316 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X1612 a_25137_864 a_23136_447 a_24913_864 VDD.t1894 pfet_06v0 ad=0.1826p pd=1.71u as=0.1079p ps=0.935u w=0.415u l=0.5u
X1613 VSS.t312 a_21772_n11428.t10 a_13623_n14874.t5 VSS.t311 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1614 a_34576_1204 a_32108_n2332.t20 VSS.t4201 VSS.t4200 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1615 VDD.t3625 a_34649_n2412 a_25836_n1236.t7 VDD.t3624 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1616 a_13623_n14874.t4 a_21772_n11428.t11 VSS.t314 VSS.t313 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1617 VDD.t373 a_10778_2852.t22 a_10712_4516.t26 VDD.t372 pfet_03v3 ad=1.82p pd=6.9u as=0.728p ps=3.32u w=2.8u l=0.28u
X1618 a_25020_n11383 a_22140_n6694.t8 a_35120_n9412 VDD.t4061 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X1619 a_32533_n12376 a_32413_n12996 a_31789_n12996 VDD.t877 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1620 a_38380_n17349 a_38292_n17252 VSS.t2771 VSS.t2770 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1621 VDD.t1338 a_29420_n17349 a_29332_n17252 VDD.t1337 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1622 a_n263_3472.t5 a_22444_2253.t14 VSS.t2427 VSS.t2426 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1623 a_46108_n4372 a_46020_n4328 VSS.t3648 VSS.t3647 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1624 a_34089_n10252 a_24481_761.t41 VDD.t730 VDD.t729 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X1625 VDD.t4113 a_25940_n17606.t6 a_21772_n12996 VDD.t4112 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1626 a_38380_n14213 a_38292_n14116 VSS.t3673 VSS.t3672 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1627 VDD.t3839 a_41852_n12212 a_41764_n12168 VDD.t3838 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1628 a_36140_n17349 a_36052_n17252 VSS.t2974 VSS.t2973 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1629 a_32412_n13648 a_31960_n13648 VDD.t3527 VDD.t3526 pfet_06v0 ad=0.2028p pd=1.3u as=0.45p ps=2.02u w=0.78u l=0.5u
X1630 a_33216_1944.t2 a_25084_1564 VSS.t1174 VSS.t1173 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1631 a_33416_n4240 a_33015_n4284 a_32359_n4372 VSS.t2879 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1632 a_27134_n9816 a_26470_n9322 VSS.t3213 VSS.t3212 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1633 a_27952_n14432 a_27804_n14165 a_27784_n14432 VSS.t1408 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1634 VSS.t1796 a_25539_n407.t3 a_25759_1944 VSS.t1795 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X1635 a_11087_n7460.t18 a_11023_n6840.t26 VSS.t105 VSS.t72 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X1636 a_36140_n14213 a_36052_n14116 VSS.t2942 VSS.t2855 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1637 VDD.t1813 a_39612_n10644 a_39524_n10600 VDD.t1812 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1638 VSS.t3705 a_34649_n2412 a_25836_n1236.t1 VSS.t3704 nfet_06v0 ad=0.2119p pd=1.335u as=0.2119p ps=1.335u w=0.815u l=0.6u
X1639 a_42300_n7508 a_42212_n7464 VSS.t3017 VSS.t3016 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1640 a_32152_n13692 a_31559_n13692 a_32888_n13248 VSS.t4074 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1641 a_27672_n3543 a_27932_n3543 VDD.t3777 VDD.t3776 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X1642 a_13501_n6460.t9 a_11023_n6840.t27 a_11087_n7460.t24 VDD.t112 pfet_03v3 ad=1.82p pd=6.9u as=0.728p ps=3.32u w=2.8u l=0.28u
X1643 a_23108_n12080 a_21940_n11684 a_22904_n12080 VDD.t2191 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1644 a_11087_n18172.t15 a_11023_n17552.t27 a_13501_n17172.t15 VDD.t404 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1645 VSS.t1880 a_30740_n7464 a_31936_n6592 VSS.t1879 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1646 a_24233_n13388 a_23816_n13248 a_24609_n13248 VSS.t4289 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X1647 a_45212_n1669 a_45124_n1572 VSS.t3294 VSS.t3293 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1648 VDD.t3829 a_24828_n18917 a_24740_n18820 VDD.t1584 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1649 a_22276_n1572.t1 a_21828_n1931 VDD.t3835 VDD.t3834 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X1650 a_11023_n6840.t7 a_13623_n6840.t27 VSS.t732 VSS.t731 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1651 a_10778_2852.t5 a_10712_4516.t39 VSS.t347 VSS.t346 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
D43 a_22444_332.t15 VDD.t2 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1652 a_27055_n12168 a_26431_n12168 a_26887_n12168 VDD.t3177 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1653 a_32108_n2332.t12 a_35456_n4628.t14 VDD.t4087 VDD.t4086 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1654 VDD.t3557 a_43756_n5940 a_43668_n5896 VDD.t3556 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1655 a_24609_n10112 a_23072_n13432.t49 VSS.t506 VSS.t505 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X1656 a_39612_n16916 a_39524_n16872 VSS.t1764 VSS.t1763 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1657 a_34953_n1572 a_34223_n1976 VSS.t2407 VSS.t2406 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X1658 a_22016_n13665 a_21604_n13252 VSS.t2218 VSS.t2217 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1659 a_34068_n4 a_33508_n408 a_33940_n408 VSS.t4323 nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X1660 VDD.t3052 a_24731_n3124.t2 a_30104_n1148 VDD.t3051 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1661 a_22016_n10529 a_21604_n10116 VSS.t3448 VSS.t3447 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1662 a_36588_n18917 a_36500_n18820 VSS.t3907 VSS.t3906 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1663 a_34367_1619 a_33467_1116 VDD.t3647 VDD.t3646 pfet_06v0 ad=0.1313p pd=1.025u as=0.29465p ps=1.74u w=0.505u l=0.5u
X1664 VSS.t1730 a_29744_n15604.t14 a_23072_n13432.t3 VSS.t1729 nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1665 VSS.t3528 a_33999_n1400 a_34475_n1976 VSS.t3527 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X1666 VDD.t3255 a_28454_n2424 a_23703_n5156.t1 VDD.t3254 pfet_06v0 ad=0.4941p pd=2.03u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1667 VDD.t1351 a_42188_n15781 a_42100_n15684 VDD.t1350 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1668 VDD.t2828 a_25577_n14956 a_25472_n14816 VDD.t2827 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X1669 a_27154_n13736 a_26470_n13736 VDD.t1210 VDD.t1209 pfet_06v0 ad=61.199993f pd=0.7u as=0.1656p ps=1.28u w=0.36u l=0.5u
X1670 a_25895_n2624 a_25547_n2445 a_24771_n2804 VSS.t3977 nfet_06v0 ad=0.1989p pd=1.465u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1671 VDD.t3940 a_45660_n7508 a_45572_n7464 VDD.t3939 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1672 VDD.t2619 a_21692_n13308.t20 a_29332_n11301 VDD.t2618 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X1673 a_23072_n13432.t4 a_29744_n15604.t15 VSS.t1732 VSS.t1731 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1674 VDD.t1938 a_42188_n12645 a_42100_n12548 VDD.t1937 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1675 a_34348_n18917 a_34260_n18820 VSS.t929 VSS.t928 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1676 VSS.t891 a_4001_4292.t8 a_10778_2852.t12 VSS.t350 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1677 VDD.t3916 a_45660_n4372 a_45572_n4328 VDD.t3915 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1678 a_24233_n10252 a_23072_n13432.t50 VDD.t502 VDD.t501 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X1679 a_43644_n18484 a_43556_n18440 VSS.t986 VSS.t985 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1680 a_46556_n13780 a_46468_n13736 VSS.t1032 VSS.t1031 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1681 a_30866_n3844 a_25836_n1236.t11 a_30662_n3844 VSS.t1105 nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1682 a_46556_n10644 a_46468_n10600 VSS.t1146 VSS.t1145 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1683 a_43644_n15348 a_43556_n15304 VSS.t1775 VSS.t1774 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1684 OUT[4].t9 a_41392_1944.t14 VDD.t1385 VDD.t1384 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1685 VDD.t2105 a_34895_376 a_35351_398 VDD.t2104 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1686 a_36408_n320 a_35568_n4 a_36120_n4 VSS.t4092 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1687 VSS.t1951 a_33832_n8572 a_25612_n6679 VSS.t1950 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X1688 a_41404_n18484 a_41316_n18440 VSS.t1388 VSS.t1387 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D44 a_23072_n13432.t51 VDD.t503 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1689 a_46668_n3237 a_46580_n3140 VSS.t3913 VSS.t3912 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1690 VDD.t2331 a_44540_n9076 a_44452_n9032 VDD.t2330 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1691 a_31459_n14564 a_31789_n14564 a_31909_n14520 VSS.t2562 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X1692 VDD.t1361 a_28492_332 a_28336_376 VDD.t1360 pfet_06v0 ad=0.4392p pd=1.94u as=0.4758p ps=2u w=1.22u l=0.5u
X1693 a_11087_n23528.t40 a_2167_3472.t62 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X1694 VDD.t2399 a_45660_n15348 a_45572_n15304 VDD.t2398 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1695 a_41404_n15348 a_41316_n15304 VSS.t2970 VSS.t2969 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1696 a_42157_n660 a_34428_n452.t3 VDD.t2973 VDD.t2972 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1697 VDD.t1057 a_21916_n6694.t7 a_29532_n4372.t0 VDD.t1056 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1698 VDD.t221 a_13623_n22908.t17 a_11023_n22908.t17 VDD.t220 pfet_03v3 ad=1.82p pd=6.9u as=0.728p ps=3.32u w=2.8u l=0.28u
X1699 VSS.t1308 a_21804_n2273.t6 a_24516_n14475 VSS.t1307 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1700 a_25795_n2716.t1 a_21692_n5468.t20 VDD.t395 VDD.t394 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X1701 VDD.t31 a_24815_n3588.t13 a_29076_n8292.t1 VDD.t30 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1702 VDD.t66 a_21772_n8292.t13 a_13623_n17552.t14 VDD.t65 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
D45 VSS.t507 a_23072_n13432.t52 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1703 VDD.t260 a_13623_n9518.t16 a_11023_n9518.t16 VDD.t259 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1704 a_27605_n9032 a_27485_n8500 a_26861_n8567 VDD.t955 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1705 a_37372_n12212 a_37284_n12168 VSS.t2903 VSS.t2902 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1706 VDD.t3237 a_44540_n15348 a_44452_n15304 VDD.t3236 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1707 a_38828_n9509 a_38740_n9412 VSS.t3966 VSS.t3965 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1708 a_32158_n12212 a_31961_n11340 VSS.t4090 VSS.t4089 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1709 a_11023_n22908.t16 a_13623_n22908.t18 VDD.t223 VDD.t222 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1710 a_30555_n2729 a_29900_n10600.t5 VDD.t3863 VDD.t3862 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1711 a_41292_n9509 a_41204_n9412 VSS.t3827 VSS.t3826 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1712 a_36252_n12212 a_36164_n12168 VSS.t3454 VSS.t3453 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1713 VDD.t2996 a_29532_n20052 a_29444_n20008 VDD.t2995 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1714 a_11087_n23528.t41 a_2167_3472.t61 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X1715 VDD.t3278 a_42300_n15348 a_42212_n15304 VDD.t3277 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1716 VDD.t2417 a_22668_n14864.t2 a_22264_n8988 VDD.t2416 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1717 VDD.t2259 a_28300_n15348 a_28437_n13705 VDD.t2258 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1718 a_43725_908 a_40260_n408 VSS.t2255 VSS.t2254 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1719 a_31235_n9860 a_31565_n9860 a_31685_n9262 VDD.t2211 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1720 VDD.t3352 a_28412_n20052 a_28324_n20008 VDD.t3351 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1721 VSS.t474 a_21772_1116.t9 a_13623_n4162.t4 VSS.t4 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1722 a_41336_n407 a_25539_n407.t4 VSS.t1798 VSS.t1797 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X1723 a_43980_n11077 a_43892_n10980 VSS.t2699 VSS.t2698 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1724 VDD.t2341 a_22444_2253.t15 a_n263_3472.t11 VDD.t2340 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1725 OUT[0].t0 a_29408_1944.t15 VSS.t3993 VSS.t3992 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1726 a_29176_n7819 a_29076_n8292.t6 a_28972_n7819 VDD.t440 pfet_06v0 ad=0.58035p pd=2.155u as=0.2847p ps=1.615u w=1.095u l=0.5u
X1727 a_28636_n16916 a_28548_n16872 VSS.t1235 VSS.t1234 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1728 OUT[5].t15 a_44640_1944.t10 VDD.t240 VDD.t239 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1729 a_27452_n2716 a_25940_n17606.t7 a_28583_n3140 VDD.t4114 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1730 VDD.t1619 a_42972_n20485 a_42884_n20388 VDD.t1618 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1731 VSS.t2756 a_11023_n4162.t26 a_2167_3472.t32 VDD.t2692 pfet_03v3 ad=0.728p pd=3.32u as=1.82p ps=6.9u w=2.8u l=0.28u
X1732 VDD.t1445 a_26531_n8639 a_22712_n7420 VDD.t1425 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1733 a_41740_n11077 a_41652_n10980 VSS.t2570 VSS.t2569 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1734 VDD.t2265 a_29980_n18484 a_29892_n18440 VDD.t2264 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1735 a_45772_n101 a_45684_n4 VSS.t3853 VSS.t3852 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1736 a_46556_n4372 a_46468_n4328 VSS.t2459 VSS.t2458 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1737 a_41740_n7941 a_41652_n7844 VSS.t1921 VSS.t1920 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1738 a_36140_n13780 a_36052_n13736 VSS.t2349 VSS.t2348 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1739 OUT[2].t9 a_37024_1944.t14 VDD.t1699 VDD.t1698 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1740 a_25076_n4.t1 a_24628_n363 VDD.t1907 VDD.t1906 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X1741 a_46108_n1236 a_46020_n1192 VSS.t2461 VSS.t2460 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1742 a_40620_n11077 a_40532_n10980 VSS.t2351 VSS.t2350 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1743 a_21692_n16916 a_21604_n16872 VSS.t1746 VSS.t1745 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1744 VSS.t401 a_21692_n5468.t21 a_22724_860.t0 VSS.t400 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1745 VDD.t2270 a_38156_n7941 a_38068_n7844 VDD.t2269 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1746 VDD.t2645 a_40732_n20485 a_40644_n20388 VDD.t2644 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1747 a_11087_n20850.t4 a_11023_n20230.t24 a_13501_n19850.t7 VDD.t1844 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1748 VSS.t2095 a_137_4292 a_3025_2852 VSS.t2094 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X1749 a_11087_n7460.t4 a_13623_n6840.t28 a_13501_n6460.t4 VSS.t733 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1750 VDD.t2646 a_34796_n13780 a_34708_n13736 VDD.t1419 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D46 a_21692_n6694.t13 VDD.t637 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1751 VDD.t2369 a_44092_n10644 a_44004_n10600 VDD.t2368 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1752 VSS.t247 a_13623_n9518.t17 a_11023_n9518.t7 VSS.t246 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1753 a_32668_n18484 a_32580_n18440 VSS.t2354 VSS.t2353 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1754 VSS.t2429 a_22444_2253.t16 a_n263_3472.t4 VSS.t2428 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1755 a_26796_1515 a_26488_1564 VSS.t2983 VSS.t2982 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X1756 a_25895_n2624 a_23072_n13432.t53 VDD.t505 VDD.t504 pfet_06v0 ad=0.1521p pd=1.105u as=0.4149p ps=2.65u w=0.585u l=0.5u
X1757 a_30555_n2729 a_22220_690.t9 VDD.t781 VDD.t780 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X1758 a_34736_n3840 a_33015_n4284 a_33608_n4284 VDD.t2813 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1759 a_11023_n9518.t6 a_13623_n9518.t18 VSS.t249 VSS.t248 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X1760 a_45660_n1669 a_45572_n1572 VSS.t3116 VSS.t1559 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1761 VDD.t2371 a_37036_n9509 a_36948_n9412 VDD.t2370 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1762 VDD.t582 a_13623_n20230.t26 a_11023_n20230.t17 VDD.t581 pfet_03v3 ad=1.82p pd=6.9u as=0.728p ps=3.32u w=2.8u l=0.28u
X1763 a_42456_1248 a_41616_1564 a_42168_1564 VSS.t2822 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1764 a_22444_332.t5 a_27259_804.t9 a_29560_n3544 VSS.t855 nfet_06v0 ad=0.4161p pd=1.905u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1765 a_11023_n20230.t16 a_13623_n20230.t27 VDD.t584 VDD.t583 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1766 a_30428_n18484 a_30340_n18440 VSS.t2467 VSS.t2466 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1767 a_30604_1515 a_30296_1564 VDD.t3561 VDD.t3560 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X1768 VDD.t2509 a_26271_n1400 a_26727_n1422 VDD.t2508 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1769 a_30676_n7844 a_30228_n8203 VSS.t3719 VSS.t3718 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X1770 a_44092_n16916 a_44004_n16872 VSS.t1853 VSS.t1852 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1771 VSS.t381 a_10778_2852.t23 a_10712_4516.t15 VSS.t380 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1772 a_11087_n18172.t32 a_2167_3472.t78 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X1773 a_29687_n13252 a_24964_n14116 VSS.t1911 VSS.t1910 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1774 VSS.t3634 a_24233_n844 a_24128_n704 VSS.t3633 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X1775 VDD.t4116 a_25940_n17606.t8 a_22444_n5156 VDD.t4115 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1776 a_47197_908 a_43644_n705 VDD.t2767 VDD.t2766 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1777 a_25412_n5895 a_21692_n6694.t14 a_25600_n5895 VDD.t638 pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1778 VSS.t61 a_11023_n14874.t27 a_11087_n15494.t26 VSS.t60 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1779 VSS.t2757 a_11023_n4162.t27 VSS.t2757 VSS.t62 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.28u
X1780 a_38828_n11077 a_38740_n10980 VSS.t2360 VSS.t2359 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1781 VDD.t2511 a_29196_n18917 a_29108_n18820 VDD.t2510 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1782 a_21812_n6643 a_21692_n6694.t15 VSS.t683 VSS.t682 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X1783 a_32309_n9816 a_32189_n9860 a_31565_n9860 VSS.t2715 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X1784 a_32732_n10556 a_32424_n10512 VSS.t4254 VSS.t4253 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X1785 a_24760_n11383 a_25020_n11383 VDD.t1288 VDD.t1287 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X1786 a_11087_n18172.t33 a_2167_3472.t77 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X1787 VSS.t359 a_26440_n5940.t8 a_21692_n5468.t6 VSS.t358 nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
D47 a_24481_761.t42 VDD.t731 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1788 VDD.t1059 a_21916_n6694.t8 a_28736_n4633.t4 VDD.t1058 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X1789 VDD.t3984 a_29532_n10311 a_29444_n10116 VDD.t3983 pfet_06v0 ad=0.35315p pd=1.96u as=0.2486p ps=2.01u w=0.565u l=0.5u
X1790 VDD.t2379 a_31996_n20485 a_31908_n20388 VDD.t2378 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1791 VDD.t4052 a_22140_n16916 a_22052_n16872 VDD.t4051 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1792 VDD.t4054 a_42188_n7941 a_42100_n7844 VDD.t4053 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1793 a_24220_n15260 a_23912_n15216 VDD.t938 VDD.t937 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X1794 a_47900_n1236 a_47812_n1192 VSS.t1182 VSS.t1181 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1795 a_33868_n4240 a_33416_n4240 VDD.t3093 VDD.t35 pfet_06v0 ad=0.2028p pd=1.3u as=0.45p ps=2.02u w=0.78u l=0.5u
X1796 VDD.t1432 a_42188_n4805 a_42100_n4708 VDD.t1431 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1797 VSS.t2093 a_137_4292 a_4001_4292.t2 VSS.t2092 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X1798 a_32340_n5112 a_30555_n2729 VSS.t3056 VSS.t3055 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1799 VSS.t106 a_11023_n6840.t28 a_11087_n7460.t17 VSS.t54 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1800 a_11087_n18172.t34 a_2167_3472.t76 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X1801 VSS.t1536 a_30808_n6334 a_30616_n6221 VSS.t1535 nfet_06v0 ad=0.2016p pd=1.48u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1802 a_24380_n20052 a_24292_n20008 VSS.t4132 VSS.t3289 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1803 VDD.t4077 a_45772_n15781 a_45684_n15684 VDD.t4076 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1804 a_31656_n704 a_29444_n708 a_30716_n1148 VDD.t2745 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X1805 VDD.t72 a_21772_n8292.t14 a_13623_n17552.t13 VDD.t71 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1806 VSS.t119 a_11023_n12196.t27 a_11087_n12816.t6 VSS.t60 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1807 VDD.t899 a_45772_n12645 a_45684_n12548 VDD.t898 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1808 a_37932_n18917 a_37844_n18820 VSS.t1496 VSS.t1495 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1809 VDD.t2419 a_42636_n6373 a_42548_n6276 VDD.t2418 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1810 VDD.t1285 a_32560_n7020 a_32455_n7420 VDD.t1284 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X1811 a_22140_n20052 a_22052_n20008 VSS.t4155 VSS.t2193 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1812 VDD.t4025 a_31324_n4372 a_32132_2428 VDD.t4024 pfet_06v0 ad=0.35315p pd=1.96u as=0.2486p ps=2.01u w=0.565u l=0.5u
X1813 VDD.t4102 a_43532_n15781 a_43444_n15684 VDD.t4101 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1814 VDD.t3514 a_42636_n3237 a_42548_n3140 VDD.t3513 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1815 a_41404_n4372 a_41316_n4328 VSS.t1163 VSS.t1162 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1816 VDD.t2567 a_24573_n6724 a_24693_n6104 VDD.t2566 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1817 VDD.t2421 a_43532_n12645 a_43444_n12548 VDD.t2420 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1818 a_24481_761.t3 a_30192_n15304.t12 VDD.t2288 VDD.t1650 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1819 a_10712_4516.t25 a_10778_2852.t24 VDD.t375 VDD.t374 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1820 VSS.t964 a_39544_420 a_39352_464 VSS.t963 nfet_06v0 ad=0.2016p pd=1.48u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1821 a_32085_n7672 a_31965_n8292 a_31341_n8292 VDD.t1556 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1822 VSS.t3341 a_28454_n2424 a_23703_n5156.t0 VSS.t3340 nfet_06v0 ad=0.2911p pd=1.53u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1823 a_31628_n5940.t9 a_33496_n6659.t17 VSS.t154 VSS.t153 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X1824 a_43084_n6373 a_42996_n6276 VSS.t3218 VSS.t3217 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1825 a_47900_n13780 a_47812_n13736 VSS.t1591 VSS.t1590 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D48 a_23072_n13432.t54 VDD.t506 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1826 a_47900_n10644 a_47812_n10600 VSS.t3818 VSS.t3817 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1827 VDD.t4144 a_39164_n18484 a_39076_n18440 VDD.t4143 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1828 VDD.t855 a_21772_n3588.t10 a_13623_n20230.t12 VDD.t854 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1829 a_46668_n15781 a_46580_n15684 VSS.t3390 VSS.t3389 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1830 VDD.t903 a_30604_1515 a_30500_1564 VDD.t902 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1831 VDD.t1076 a_25836_n1236.t12 a_28736_n4633.t7 VDD.t1075 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X1832 a_38853_n5321 a_38733_n5431 VSS.t2245 VSS.t2244 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X1833 a_11023_n14874.t7 a_13623_n14874.t26 VSS.t1356 VSS.t1355 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1834 a_33653_376 a_33533_908 a_32909_841 VDD.t3053 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1835 VSS.t1924 a_11023_n20230.t25 a_11087_n20850.t5 VSS.t64 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X1836 VSS.t1358 a_13623_n14874.t27 a_11023_n14874.t8 VSS.t1357 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1837 a_39868_n408 a_29900_760.t8 a_39556_n4 VSS.t2295 nfet_06v0 ad=98.399994f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1838 a_22876_n10556 a_22568_n10512 VSS.t1133 VSS.t1132 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X1839 a_13623_n9518.t2 a_21772_n17700.t10 VDD.t1005 VDD.t1004 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1840 a_44428_n15781 a_44340_n15684 VSS.t3964 VSS.t3963 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1841 a_26553_377.t1 a_25817_804 VDD.t3141 VDD.t3140 pfet_06v0 ad=0.6561p pd=3.51u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1842 a_36744_n1954 a_36388_n1572 VSS.t1071 VSS.t1070 nfet_06v0 ad=0.1584p pd=1.6u as=0.151p ps=1.185u w=0.36u l=0.6u
X1843 a_11087_n20850.t6 a_11023_n20230.t26 VSS.t1925 VSS.t66 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1844 a_13623_n12196.t15 a_21772_n14564.t6 VDD.t2002 VDD.t2001 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1845 a_13623_n4162.t3 a_21772_1116.t10 VSS.t662 VSS.t661 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1846 a_37844_1564 a_37396_1205 VSS.t2846 VSS.t2845 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X1847 a_22444_2253.t5 a_24236_2258.t5 VDD.t2348 VDD.t2347 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1848 VDD.t3676 a_30900_n9032 a_21692_n6694.t1 VDD.t3675 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
D49 a_21692_n6694.t16 VDD.t639 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1849 a_11023_n17552.t5 a_13623_n17552.t26 VSS.t86 VSS.t85 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1850 VDD.t242 a_44640_1944.t11 OUT[5].t14 VDD.t241 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
D50 VSS.t792 a_24481_761.t43 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1851 a_39056_820 a_32108_n2332.t21 VSS.t4203 VSS.t4202 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1852 a_34708_n5896.t5 a_33776_n5896.t12 VSS.t876 VSS.t875 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1853 a_26983_n12728 a_27744_n12908 a_27535_n12493 VSS.t1569 nfet_06v0 ad=0.2007p pd=1.475u as=94.5f ps=0.885u w=0.36u l=0.6u
X1854 VSS.t195 a_11023_n22908.t26 a_11087_n23528.t26 VSS.t70 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1855 a_11087_n23528.t25 a_11023_n22908.t27 VSS.t196 VSS.t72 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X1856 a_n263_3472.t3 a_22444_2253.t17 VSS.t2431 VSS.t2430 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1857 VDD.t2810 a_37484_n9509 a_37396_n9412 VDD.t2809 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D51 VSS.t684 a_21692_n6694.t17 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1858 a_11087_n20850.t33 a_2167_3472.t20 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X1859 a_25636_n14520 a_21996_n12996.t7 a_24965_n9860 VSS.t3573 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1860 a_33216_1944.t1 a_25084_1564 VSS.t1172 VSS.t1171 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1861 VDD.t2365 a_46108_n1236 a_46020_n1192 VDD.t2194 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1862 a_35456_n4628.t1 a_34708_n5896.t21 VSS.t862 VSS.t861 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1863 a_31548_n10172.t4 a_33496_n8222.t12 VSS.t298 VSS.t297 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1864 a_11023_n12196.t7 a_13623_n12196.t26 VSS.t1832 VSS.t1831 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1865 VDD.t1839 a_34796_n15781 a_34708_n15684 VDD.t1201 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1866 VDD.t556 a_13623_n4162.t23 a_11023_n4162.t17 VDD.t555 pfet_03v3 ad=1.82p pd=6.9u as=0.728p ps=3.32u w=2.8u l=0.28u
X1867 VSS.t1834 a_13623_n12196.t27 a_11023_n12196.t8 VSS.t1833 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1868 a_29744_1564 a_29332_1243 VDD.t2515 VDD.t2514 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
D52 a_24481_761.t44 VDD.t732 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1869 a_26956_n18917 a_26868_n18820 VSS.t966 VSS.t965 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1870 a_13501_n14494.t3 a_13623_n14874.t28 a_11087_n15494.t3 VSS.t1359 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X1871 a_35849_n1192 a_35119_n1170 VDD.t2863 VDD.t2862 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X1872 VDD.t1924 a_40060_n4805 a_39972_n4708 VDD.t1546 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1873 a_13623_n17552.t3 a_21772_n8292.t15 VSS.t427 VSS.t426 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1874 a_24069_n9816 a_23949_n9860 VSS.t2004 VSS.t2003 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X1875 a_47900_n5940 a_47812_n5896 VSS.t3871 VSS.t3870 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1876 a_29211_n6724 a_29559_n6456 VDD.t2907 VDD.t2906 pfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X1877 a_32543_n9032 a_31919_n9032 a_32375_n9032 VDD.t2144 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1878 VDD.t913 a_46220_n101 a_46132_n4 VDD.t912 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1879 VDD.t290 a_33496_n8222.t13 a_31548_n10172.t13 VDD.t289 pfet_06v0 ad=0.367p pd=1.92u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1880 VDD.t1727 a_31664_n13292 a_31559_n13692 VDD.t1726 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X1881 VDD.t2431 a_35849_n1192 a_36192_1248 VDD.t2430 pfet_06v0 ad=0.3432p pd=2.44u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1882 VSS.t4148 a_23619_n9860 a_22264_n10556 VSS.t4147 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1883 a_42188_n11077 a_42100_n10980 VSS.t4173 VSS.t4172 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1884 a_25620_n5412 a_24672_n11339 VSS.t1968 VSS.t1967 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1885 a_21772_n20836.t2 a_23564_n20836 VSS.t944 VSS.t943 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1886 a_30296_1564 a_29744_1564 a_30092_1564 VDD.t1112 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1887 VSS.t701 a_21772_n20836.t14 a_13623_n6840.t3 VSS.t700 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1888 a_34895_n1192 a_34271_n1192 a_34727_n1192 VDD.t1349 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1889 VDD.t164 a_33496_n6659.t18 a_31628_n5940.t28 VDD.t163 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1890 VDD.t3233 a_23619_n12996 a_22264_n13692 VDD.t3232 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1891 VSS.t4266 a_37844_1564 a_38256_1564.t3 VSS.t4265 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1892 VSS.t2710 a_47197_908 a_47317_952 VSS.t2709 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1893 a_13501_n11816.t13 a_13623_n12196.t28 a_11087_n12816.t23 VSS.t1835 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X1894 a_22544_n4690 a_22444_n5156 VDD.t2519 VDD.t2518 pfet_06v0 ad=0.4248p pd=1.94u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1895 a_47116_n18917 a_47028_n18820 VSS.t1974 VSS.t1973 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1896 a_13501_n17172.t6 a_13623_n17552.t27 a_11087_n18172.t6 VSS.t87 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1897 VDD.t734 a_24481_761.t45 a_24041_816 VDD.t733 pfet_06v0 ad=0.4149p pd=2.65u as=0.1521p ps=1.105u w=0.585u l=0.5u
X1898 VDD.t4136 a_41292_n1669 a_41204_n1572 VDD.t4135 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1899 VSS.t794 a_24481_761.t46 a_33955_1240 VSS.t793 nfet_06v0 ad=0.1224p pd=1.04u as=0.134p ps=1.1u w=0.36u l=0.6u
X1900 a_41292_n18917 a_41204_n18820 VSS.t1184 VSS.t1183 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1901 a_41852_n4372 a_41764_n4328 VSS.t1613 VSS.t1612 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1902 a_30348_n6980 a_28736_n4633.t21 a_30036_n7464 VSS.t1072 nfet_06v0 ad=98.399994f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1903 VDD.t4138 a_22140_n15781 a_22052_n15684 VDD.t1218 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1904 a_37947_332 a_38295_332 VDD.t1182 VDD.t1181 pfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X1905 a_21772_n11428.t2 a_23564_n11428 VSS.t1752 VSS.t1751 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1906 a_40172_n18917 a_40084_n18820 VSS.t1186 VSS.t1185 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1907 VSS.t316 a_21772_n11428.t12 a_13623_n14874.t3 VSS.t315 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1908 a_33308_n7376 a_32856_n7376 VDD.t2752 VDD.t2751 pfet_06v0 ad=0.2028p pd=1.3u as=0.45p ps=2.02u w=0.78u l=0.5u
X1909 VDD.t2838 a_28300_n18917 a_28212_n18820 VDD.t2837 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D53 VSS.t1899 CLK.t6 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1910 VDD.t2844 a_43644_n12212 a_43556_n12168 VDD.t2843 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1911 a_24684_n16432 a_25831_n11428 a_25767_n11383 VSS.t1859 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1912 VSS.t3323 a_29263_n3588.t2 a_29199_n3543 VSS.t3322 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1913 a_32189_n9860 a_32581_n9860 VSS.t2905 VSS.t2904 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1914 VDD.t3239 a_41404_n12212 a_41316_n12168 VDD.t3238 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1915 a_43833_1204 a_43416_1248 a_44209_1248 VSS.t1650 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X1916 VDD.t3155 a_43532_n9509 a_43444_n9412 VDD.t3154 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1917 a_11087_n23528.t10 a_11023_n22908.t28 a_13501_n22528.t16 VDD.t209 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1918 VDD.t1078 a_25836_n1236.t13 a_29956_n2760 VDD.t1077 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1919 a_13501_n19850.t15 a_13623_n20230.t28 a_11087_n20850.t25 VSS.t625 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1920 a_26531_n10207 a_26861_n10135 a_26981_n10578 VDD.t1543 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1921 VDD.t2439 a_38312_n1975 a_32636_n2020 VDD.t2438 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1922 a_39477_n5320 a_39357_n5364 a_38733_n5431 VSS.t1193 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X1923 a_39948_n7941 a_39860_n7844 VSS.t2897 VSS.t2896 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1924 a_11087_n20850.t32 a_2167_3472.t18 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X1925 a_23036_n15781 a_22948_n15684 VSS.t1872 VSS.t1871 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1926 VSS.t476 a_21772_1116.t11 a_13623_n4162.t2 VSS.t475 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1927 a_13623_n20230.t11 a_21772_n3588.t11 VDD.t857 VDD.t856 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1928 a_34000_n3140 a_33588_n3461 VDD.t3340 VDD.t3339 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X1929 VDD.t2929 a_26643_n8292 a_23887_n5156 VDD.t2928 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1930 VSS.t1059 a_24233_n8684 a_24128_n8544 VSS.t1058 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X1931 VSS.t3691 a_31961_1204 a_31856_1248 VSS.t3690 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X1932 VDD.t3122 a_35288_n1975 a_34248_n3310 VDD.t3121 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1933 a_34708_n5896.t4 a_33776_n5896.t13 VSS.t878 VSS.t877 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1934 OUT[5].t13 a_44640_1944.t12 VDD.t244 VDD.t243 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1935 VSS.t3031 a_24233_n5548 a_24128_n5408 VSS.t3030 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X1936 a_26796_1515 a_26488_1564 VDD.t2911 VDD.t2910 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
D54 VSS.t795 a_24481_761.t47 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1937 a_46556_n1236 a_46468_n1192 VSS.t3611 VSS.t3610 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1938 VDD.t2594 a_26047_n4328 a_26503_n4306 VDD.t2593 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1939 a_11087_n20850.t34 a_2167_3472.t21 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X1940 a_26098_n13736 a_25642_n13736 VDD.t1185 VDD.t1184 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1941 a_10712_4516.t14 a_10778_2852.t25 VSS.t383 VSS.t382 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1942 a_34460_n16916 a_34372_n16872 VSS.t3441 VSS.t3440 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1943 VDD.t3717 a_25132_n16432 a_23608_n15260 VDD.t3716 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1944 a_22444_332.t1 a_29920_n3900.t15 VDD.t610 VDD.t609 pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X1945 a_27205_n15534 a_27085_n16132 VDD.t1882 VDD.t1881 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X1946 VDD.t1159 a_46556_n1236 a_46468_n1192 VDD.t1158 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1947 a_39804_464 a_39352_464 VDD.t3219 VDD.t3218 pfet_06v0 ad=0.2028p pd=1.3u as=0.45p ps=2.02u w=0.78u l=0.5u
X1948 a_32220_n16916 a_32132_n16872 VSS.t2598 VSS.t2597 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1949 a_21772_n8292.t3 a_23564_n8292 VSS.t1223 VSS.t1222 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1950 a_24128_n10112 a_21604_n10116 a_23816_n10112 VSS.t3446 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1951 a_11087_n23528.t6 a_13623_n22908.t19 a_13501_n22528.t6 VSS.t213 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1952 a_47116_n101 a_47028_n4 VSS.t1633 VSS.t1632 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1953 VDD.t2445 a_38716_n7508 a_38628_n7464 VDD.t2444 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1954 a_46556_n18484 a_46468_n18440 VSS.t1213 VSS.t1212 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1955 a_24116_n15216 a_23072_n13432.t55 VDD.t508 VDD.t507 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X1956 VSS.t3846 a_21692_2431 a_21604_2475 VSS.t3845 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1957 VSS.t2433 a_22444_2253.t18 a_n263_3472.t2 VSS.t2432 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1958 VDD.t1007 a_21772_n17700.t11 a_13623_n9518.t2 VDD.t1006 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1959 a_46556_n15348 a_46468_n15304 VSS.t2972 VSS.t2971 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1960 VDD.t1579 a_32413_n14564 a_32533_n13944 VDD.t1578 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1961 VDD.t2658 a_47900_n1669 a_47812_n1572 VDD.t2657 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1962 VSS.t300 a_33496_n8222.t14 a_31548_n10172.t3 VSS.t299 nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
D55 VSS.t508 a_23072_n13432.t56 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1963 VSS.t455 a_3935_4156.t6 a_10712_4516.t3 VSS.t384 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1964 VDD.t2506 a_26796_1515 a_26692_1564 VDD.t2505 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1965 a_28076_n17349 a_27988_n17252 VSS.t3806 VSS.t1489 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1966 VDD.t2004 a_21772_n14564.t7 a_13623_n12196.t14 VDD.t2003 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1967 VSS.t439 a_33216_1944.t14 OUT[1].t6 VSS.t438 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1968 a_25524_n708 a_25836_n1236.t14 a_23404_816 VSS.t1106 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1969 a_29800_n5940.t4 a_31628_n5940.t36 VDD.t144 VDD.t143 pfet_06v0 ad=0.2952p pd=1.54u as=0.367p ps=1.92u w=0.82u l=0.5u
X1970 VDD.t2280 a_21812_n6643 a_25412_n8501 VDD.t2279 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1971 a_46108_n13780 a_46020_n13736 VSS.t2623 VSS.t2622 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1972 a_32073_n844 a_23072_n13432.t57 VDD.t510 VDD.t509 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X1973 VDD.t1555 a_31965_n8292 a_32085_n7672 VDD.t1554 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1974 VDD.t2662 a_47452_n15348 a_47364_n15304 VDD.t2661 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1975 a_24681_n7116 a_24264_n6976 a_25057_n6976 VSS.t2476 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X1976 a_46108_n10644 a_46020_n10600 VSS.t1649 VSS.t1648 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1977 VSS.t510 a_23072_n13432.t58 a_23360_n11680 VSS.t509 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1978 a_31412_n2276 a_31292_n2804 VSS.t2976 VSS.t2975 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1979 a_42188_n3237 a_42100_n3140 VSS.t1225 VSS.t1224 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1980 VSS.t2679 a_21692_n13308.t21 a_29332_n11301 VSS.t2678 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1981 VDD.t166 a_33496_n6659.t19 a_31628_n5940.t27 VDD.t165 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1982 VDD.t1258 a_24752_n8292 a_22140_n6694.t1 VDD.t1257 pfet_06v0 ad=0.35315p pd=1.96u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1983 VDD.t2300 a_40060_n9076 a_39972_n9032 VDD.t2299 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1984 VDD.t1748 a_13623_n12196.t29 a_11023_n12196.t9 VDD.t1747 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1985 a_39164_n12212 a_39076_n12168 VSS.t2390 VSS.t2389 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1986 a_45660_332 a_45572_376 VSS.t2723 VSS.t2722 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1987 a_42244_n1572 a_41684_n1976 a_42116_n1976 VSS.t2477 nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X1988 a_11023_n17552.t16 a_13623_n17552.t28 VDD.t94 VDD.t93 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1989 VDD.t2304 a_45212_n15348 a_45124_n15304 VDD.t2303 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1990 VSS.t2343 a_46243_769 a_42604_n2020 VSS.t2342 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1991 a_24128_n3840 a_21604_n3844 a_23816_n3840 VSS.t1806 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1992 VDD.t1829 a_37785_n364 a_37680_n320 VDD.t1828 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X1993 a_28791_n3543 a_25940_n17606.t9 VSS.t4183 VSS.t4182 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1994 a_31939_n6976 a_31799_n7508 a_31451_n7508 VSS.t1627 nfet_06v0 ad=0.134p pd=1.1u as=0.176p ps=1.68u w=0.4u l=0.6u
X1995 a_32413_n12996 a_28927_n10160 VSS.t2397 VSS.t2396 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1996 VSS.t1316 a_44509_n452 a_44629_n408 VSS.t1315 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1997 a_45772_n11077 a_45684_n10980 VSS.t2729 VSS.t2728 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1998 VDD.t2386 a_33900_n15781 a_33812_n15684 VDD.t2385 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1999 a_46243_769 a_46573_841 a_46693_398 VDD.t2733 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2000 a_25895_n2624 a_25795_n2716.t2 a_24771_n2804 VDD.t2355 pfet_06v0 ad=0.27805p pd=2.17u as=0.1079p ps=0.935u w=0.415u l=0.5u
X2001 a_27717_n7672 a_27597_n8292 a_26973_n8292 VDD.t2879 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2002 VDD.t4075 a_24380_n20052 a_24292_n20008 VDD.t4074 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2003 VDD.t2388 a_45884_n20485 a_45796_n20388 VDD.t2387 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2004 a_1955_4292.t0 a_n263_3472.t17 VDD.t2010 VDD.t2009 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X2005 VDD.t2024 a_48012_332 a_47924_376 VDD.t2023 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2006 VDD.t2570 a_43868_n2804 a_43780_n2760 VDD.t2569 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2007 a_22876_n4284 a_22568_n4240 VSS.t3046 VSS.t3045 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X2008 a_43532_n11077 a_43444_n10980 VSS.t2731 VSS.t2730 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D56 a_24481_761.t48 VDD.t735 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2009 a_25237_n5895 a_24233_n5548 VSS.t3029 VSS.t3028 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2010 VDD.t4100 a_22140_n20052 a_22052_n20008 VDD.t4099 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2011 a_36140_n15348 a_36052_n15304 VSS.t2856 VSS.t2855 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2012 VDD.t2578 a_41203_n799 a_39308_n452 VDD.t2577 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2013 a_21872_n9394 a_21772_n9860 VDD.t2741 VDD.t2740 pfet_06v0 ad=0.4248p pd=1.94u as=0.4972p ps=3.14u w=1.13u l=0.5u
X2014 a_23484_n16916 a_23396_n16872 VSS.t3041 VSS.t3040 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2015 VDD.t1567 a_34576_1204 a_34471_1575 VDD.t1566 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2016 a_28624_n9394 a_28519_n10160.t7 a_28644_n9815 VSS.t844 nfet_06v0 ad=0.4137p pd=1.9u as=0.2119p ps=1.335u w=0.815u l=0.6u
D57 a_22444_332.t16 VDD.t3 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2017 VDD.t2318 a_42524_n20485 a_42436_n20388 VDD.t2317 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2018 VDD.t2572 a_29532_n18484 a_29444_n18440 VDD.t2571 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2019 VDD.t2322 a_42748_n7508 a_42660_n7464 VDD.t2321 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2020 VDD.t2674 a_42748_n4372 a_42660_n4328 VDD.t2673 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2021 a_11023_n14874.t9 a_13623_n14874.t29 VDD.t1308 VDD.t1307 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2022 VDD.t2324 a_36588_n13780 a_36500_n13736 VDD.t2323 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2023 VDD.t2676 a_43980_n9509 a_43892_n9412 VDD.t2675 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2024 VDD.t2848 a_33900_n11428 a_32581_n9860 VDD.t2847 pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X2025 VDD.t2855 a_27055_n12168 a_27511_n12146 VDD.t2854 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2026 VSS.t3163 a_30451_n452 a_28456_n364 VSS.t3162 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2027 a_23619_n9860 a_23949_n9860 a_24069_n9816 VSS.t2002 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X2028 a_30903_n13780 a_31664_n13292 a_31455_n13648 VSS.t1812 nfet_06v0 ad=0.2007p pd=1.475u as=94.5f ps=0.885u w=0.36u l=0.6u
X2029 VSS.t456 a_3935_4156.t7 a_10712_4516.t4 VSS.t386 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2030 a_21772_n3588.t1 a_23564_n3588.t3 VDD.t2915 VDD.t2914 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2031 VSS.t2415 a_37452_n3888 a_32860_n2020 VSS.t2414 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X2032 a_42524_n2804 a_42436_n2760 VSS.t2739 VSS.t2738 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2033 VDD.t2396 a_45324_n6373 a_45236_n6276 VDD.t2395 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2034 VSS.t3271 a_32650_n12168 a_33126_n11592 VSS.t3270 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2035 VDD.t2682 a_45324_n3237 a_45236_n3140 VDD.t2681 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2036 VDD.t2975 a_34428_n452.t4 a_37396_1205 VDD.t2974 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X2037 a_39760_n4 a_38996_n408 a_39556_n4 VDD.t2397 pfet_06v0 ad=0.4758p pd=2u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2038 VSS.t6 a_22444_332.t17 a_36155_n10116 VSS.t5 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2039 a_35800_1248 a_34872_1619 a_35632_1248 VSS.t1466 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2040 VSS.t880 a_33776_n5896.t14 a_34708_n5896.t3 VSS.t879 nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2041 a_27884_332.t1 a_29519_n1976 VDD.t2329 VDD.t2328 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X2042 VDD.t3841 a_24771_n2804 a_24403_n2414 VDD.t3840 pfet_06v0 ad=0.3276p pd=1.62u as=0.3432p ps=2.44u w=0.78u l=0.5u
X2043 VSS.t4103 a_31324_n4372 a_32132_2428 VSS.t4102 nfet_06v0 ad=0.2344p pd=1.56u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2044 a_21772_1116.t1 a_23564_1116.t4 VSS.t3493 VSS.t3492 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2045 a_11087_n7460.t23 a_11023_n6840.t29 a_13501_n6460.t6 VDD.t113 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2046 a_30740_n7464 a_30036_n7464 VSS.t3141 VSS.t3140 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2047 a_34736_n3840 a_33120_n3884 a_33608_n4284 VSS.t3643 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2048 VDD.t246 a_44640_1944.t13 OUT[5].t12 VDD.t245 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2049 VDD.t3786 a_29800_n9815 a_22220_n12996 VDD.t1056 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2050 a_26118_n9816 a_25642_n9816 VSS.t2311 VSS.t2310 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2051 a_33364_n11384 a_29444_n4328.t7 a_32581_n9860 VSS.t1561 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2052 a_24094_n1400 a_23954_n2020 VDD.t2200 VDD.t2199 pfet_06v0 ad=61.199993f pd=0.7u as=0.1656p ps=1.28u w=0.36u l=0.5u
X2053 a_13623_n22908.t1 a_21772_n452.t9 VDD.t1596 VDD.t779 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2054 VSS.t2297 a_29900_760.t9 a_33508_n408 VSS.t2296 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2055 OUT[2].t7 a_37024_1944.t15 VSS.t1777 VSS.t1776 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2056 VDD.t4034 a_38268_n4805 a_38180_n4708 VDD.t4033 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2057 VSS.t2162 a_32158_n12212 a_32026_n12168 VSS.t2161 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X2058 VSS.t3591 a_27709_n16132 a_27829_n16088 VSS.t3590 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2059 a_25953_n14816 a_23072_n13432.t59 VSS.t512 VSS.t511 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X2060 VDD.t4265 a_31548_n20485 a_31460_n20388 VDD.t4264 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2061 a_24731_n3124.t1 a_25019_n3588.t4 a_24935_n3544 VSS.t3474 nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X2062 VSS.t1701 a_26383_n2968 a_26859_n3544 VSS.t1700 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X2063 a_26172_n20052 a_26084_n20008 VSS.t3123 VSS.t3122 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D58 VSS.t685 a_21692_n6694.t18 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2064 VDD.t2909 a_24041_816 a_23981_464 VDD.t2908 pfet_06v0 ad=0.3975p pd=2.185u as=0.101p ps=0.905u w=0.505u l=0.5u
D59 VSS.t7 a_22444_332.t18 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2065 a_37372_n5940 a_37284_n5896 VSS.t3825 VSS.t3824 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D60 a_26388_n17606.t6 VDD.t323 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2066 a_13501_n19850.t6 a_11023_n20230.t27 a_11087_n20850.t7 VDD.t1845 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2067 VDD.t2210 a_47564_n15781 a_47476_n15684 VDD.t2209 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2068 a_39724_n18917 a_39636_n18820 VSS.t2294 VSS.t2293 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2069 a_22444_2253.t2 a_24236_2258.t6 VSS.t2439 VSS.t2438 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2070 a_30576_376 a_29812_860 a_30372_376 VDD.t3504 pfet_06v0 ad=0.4758p pd=2u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2071 VSS.t2499 a_23999_n2320.t4 a_23935_n2276 VSS.t2498 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2072 a_33188_n2672 a_32020_n2276 a_32984_n2672 VDD.t3023 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2073 a_24576_n6976 a_22052_n6980 a_24264_n6976 VSS.t1554 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2074 a_28972_n8247 a_29123_n6679 a_28764_n8247 VSS.t2601 nfet_06v0 ad=0.2119p pd=1.335u as=0.4137p ps=1.9u w=0.815u l=0.6u
X2075 VDD.t4208 a_47564_n12645 a_47476_n12548 VDD.t4207 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2076 a_11087_n20850.t8 a_11023_n20230.t28 a_13501_n19850.t5 VDD.t1846 pfet_03v3 ad=0.728p pd=3.32u as=1.82p ps=6.9u w=2.8u l=0.28u
X2077 a_29846_n3844 a_25836_n1236.t15 a_29652_n3844 VSS.t1107 nfet_06v0 ad=0.1517p pd=1.19u as=0.1517p ps=1.19u w=0.82u l=0.6u
X2078 VDD.t2449 a_45324_n15781 a_45236_n15684 VDD.t2448 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2079 VDD.t2977 a_34428_n452.t5 a_34272_n4 VDD.t2976 pfet_06v0 ad=0.4392p pd=1.94u as=0.4758p ps=2u w=1.22u l=0.5u
X2080 VDD.t4214 a_45324_n12645 a_45236_n12548 VDD.t4213 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2081 a_32780_n18917 a_32692_n18820 VSS.t2549 VSS.t2548 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2082 a_30759_n2276 a_21916_n6694.t9 a_30575_n2276 VSS.t1091 nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2083 a_33496_n8222.t2 a_34708_n5896.t22 VSS.t864 VSS.t863 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2084 VSS.t251 a_13623_n9518.t19 a_11023_n9518.t5 VSS.t250 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2085 a_47900_n18484 a_47812_n18440 VSS.t1530 VSS.t1529 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2086 a_24698_n1976 a_24578_n2020 a_23954_n2020 VSS.t4294 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X2087 a_30540_n18917 a_30452_n18820 VSS.t2553 VSS.t2552 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2088 a_47900_n15348 a_47812_n15304 VSS.t2895 VSS.t2894 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2089 VDD.t2451 a_38380_n11077 a_38292_n10980 VDD.t2450 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2090 a_29420_n17349 a_29332_n17252 VSS.t993 VSS.t992 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2091 a_24481_761.t0 a_30192_n15304.t13 VDD.t2289 VDD.t1636 pfet_06v0 ad=0.4392p pd=1.94u as=0.367p ps=1.92u w=1.22u l=0.5u
X2092 VSS.t2991 a_23564_n3588.t4 a_21772_n3588.t0 VSS.t2990 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2093 a_11023_n9518.t15 a_13623_n9518.t20 VDD.t262 VDD.t261 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2094 a_41392_1944.t4 a_40196_1944 VDD.t3058 VDD.t3057 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2095 a_33488_n12996 a_28927_n10160 VDD.t2314 VDD.t2313 pfet_06v0 ad=0.2486p pd=2.01u as=0.35315p ps=1.96u w=0.565u l=0.5u
D61 a_22444_332.t19 VDD.t4 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2096 VSS.t2610 a_31076_376 a_34271_n1192 VSS.t2609 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X2097 a_23816_n13248 a_22016_n13665 a_22876_n13692 VSS.t3927 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2098 a_21996_n12996.t2 a_30584_n1954 VDD.t3510 VDD.t3509 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2099 a_11087_n15494.t25 a_11023_n14874.t28 VSS.t63 VSS.t62 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2100 VSS.t578 a_13623_n4162.t24 a_11023_n4162.t6 VSS.t577 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2101 VSS.t2395 a_28927_n10160 a_28863_n10116 VSS.t2394 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2102 a_7119_4292 a_1955_4292.t3 VSS.t1399 VSS.t1398 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X2103 a_11087_n23528.t42 a_2167_3472.t60 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X2104 a_22544_n4690 a_21996_n12996.t8 a_22564_n5112 VSS.t3574 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2105 a_43532_n4805 a_43444_n4708 VSS.t2782 VSS.t2781 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2106 VDD.t2615 a_26328_n6654.t16 a_21692_n13308.t11 VDD.t2614 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2107 VSS.t413 a_11023_n17552.t28 a_11087_n18172.t26 VSS.t64 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X2108 a_26440_n5940.t0 a_28156_n6412.t21 VDD.t122 VDD.t121 pfet_06v0 ad=0.2952p pd=1.54u as=0.367p ps=1.92u w=0.82u l=0.5u
X2109 VSS.t2671 a_26328_n6654.t17 a_21692_n13308.t2 VSS.t2670 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2110 a_30599_n12167 a_31279_n11728 VDD.t2413 VDD.t2412 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2111 a_40508_n4805 a_40420_n4708 VSS.t2564 VSS.t2563 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2112 a_11087_n10138.t23 a_13623_n9518.t21 a_13501_n9138.t16 VSS.t252 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2113 a_11087_n18172.t25 a_11023_n17552.t29 VSS.t414 VSS.t66 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2114 VDD.t1208 a_46108_n5940 a_46020_n5896 VDD.t1207 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2115 a_42972_n2804 a_42884_n2760 VSS.t1661 VSS.t1660 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2116 VDD.t2484 a_45772_n6373 a_45684_n6276 VDD.t2483 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2117 a_26719_n7464 a_26095_n7464 a_26551_n7464 VDD.t1113 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2118 a_21692_n6694.t0 a_30900_n9032 VSS.t3761 VSS.t3760 nfet_06v0 ad=0.2132p pd=1.34u as=0.2911p ps=1.53u w=0.82u l=0.6u
X2119 a_44640_1944.t5 a_44004_n1192 VDD.t2498 VDD.t2497 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2120 VDD.t1215 a_46108_n2804 a_46020_n2760 VDD.t1214 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2121 VDD.t1581 a_45772_n3237 a_45684_n3140 VDD.t1580 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2122 a_44540_n4372 a_44452_n4328 VSS.t2566 VSS.t2565 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2123 VDD.t2327 a_37452_n3888 a_32860_n2020 VDD.t2326 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2124 VDD.t989 a_36588_n15781 a_36500_n15684 VDD.t988 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2125 a_30808_n10116 a_28721_n9076.t5 a_30808_n10600 VDD.t412 pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2126 a_28748_n18917 a_28660_n18820 VSS.t1534 VSS.t1533 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2127 a_45212_n1236 a_45124_n1192 VSS.t2534 VSS.t2533 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2128 a_32108_n2332.t3 a_35456_n4628.t15 VSS.t4165 VSS.t4164 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2129 a_11087_n12816.t5 a_11023_n12196.t28 VSS.t120 VSS.t62 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2130 VDD.t1480 a_35468_n12645 a_35380_n12548 VDD.t1479 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2131 VDD.t1681 a_34348_n15781 a_34260_n15684 VDD.t1328 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2132 a_26508_n18917 a_26420_n18820 VSS.t2536 VSS.t2535 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2133 a_43221_951 a_43101_841 VSS.t1928 VSS.t1927 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X2134 VDD.t3261 a_31405_n452 a_31525_168 VDD.t3260 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2135 a_46108_n9076 a_46020_n9032 VSS.t3414 VSS.t3413 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2136 VDD.t999 a_46220_n9509 a_46132_n9412 VDD.t998 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2137 VDD.t1944 a_37859_377 a_39748_2475 VDD.t1943 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X2138 a_24716_1208.t0 a_31961_1204 VSS.t3689 VSS.t3688 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
D62 a_25940_n17606.t10 VDD.t4117 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2139 a_35804_n18484 a_35716_n18440 VSS.t2017 VSS.t2016 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2140 a_38716_n13780 a_38628_n13736 VSS.t2019 VSS.t2018 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2141 VDD.t6 a_22444_332.t20 a_22340_376 VDD.t5 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2142 a_11023_n6840.t8 a_13623_n6840.t29 VDD.t672 VDD.t671 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2143 a_35120_n9412 a_28721_n9076.t6 VDD.t414 VDD.t413 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2144 VSS.t942 a_23564_n20836 a_21772_n20836.t1 VSS.t941 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2145 a_27778_n13161 a_27302_n13160 a_27526_n13714 VSS.t2537 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X2146 a_38716_n10644 a_38628_n10600 VSS.t3103 VSS.t3102 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2147 a_26907_n11592 a_26431_n12168 VSS.t3260 VSS.t3259 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2148 a_13623_n6840.t2 a_21772_n20836.t15 VSS.t668 VSS.t667 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2149 VSS.t3495 a_23564_1116.t5 a_21772_1116.t2 VSS.t3494 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2150 a_43833_1204 a_24481_761.t49 VDD.t737 VDD.t736 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X2151 a_31872_n10529 a_31460_n10116 VSS.t1323 VSS.t1322 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2152 VDD.t3014 a_37820_n15348 a_37732_n15304 VDD.t3013 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2153 VDD.t2542 a_31076_376 a_34271_n1192 VDD.t2541 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2154 a_22444_332.t4 a_27259_804.t10 a_29560_n3544 VSS.t856 nfet_06v0 ad=0.4161p pd=1.905u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2155 a_13501_n14494.t15 a_11023_n14874.t29 a_11087_n15494.t15 VDD.t77 pfet_03v3 ad=1.82p pd=6.9u as=0.728p ps=3.32u w=2.8u l=0.28u
X2156 VSS.t1926 a_11023_n20230.t29 a_11087_n20850.t9 VSS.t68 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2157 VDD.t1602 a_30732_332.t2 a_35940_2475 VDD.t1601 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X2158 a_47564_n101 a_47476_n4 VSS.t3481 VSS.t3480 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2159 a_27019_n11384 a_26543_n11384 VSS.t2022 VSS.t2021 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2160 a_27337_1944.t1 a_26607_1966 VDD.t3668 VDD.t3667 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X2161 VDD.t2081 a_32732_n10556 a_32628_n10512 VDD.t2080 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2162 a_43084_n18917 a_42996_n18820 VSS.t1247 VSS.t1246 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2163 a_23972_864 a_23136_447 a_23728_464 VSS.t1970 nfet_06v0 ad=62.1f pd=0.705u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2164 VSS.t468 a_29076_n8292.t7 a_31032_n10116 VSS.t467 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2165 VSS.t441 a_33216_1944.t15 OUT[1].t5 VSS.t440 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2166 a_23999_n2320.t0 a_24233_n844 VSS.t3632 VSS.t3631 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
D63 a_22140_n6694.t9 VDD.t4062 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2167 VDD.t1234 a_38268_n9076 a_38180_n9032 VDD.t1233 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2168 VSS.t197 a_11023_n22908.t29 a_11087_n23528.t24 VSS.t54 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2169 a_21692_n5468.t12 a_26440_n5940.t9 VDD.t348 VDD.t347 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2170 VDD.t1236 a_37708_n7941 a_37620_n7844 VDD.t1235 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2171 a_29800_n9815 a_28624_n9394 VSS.t4286 VSS.t4285 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X2172 VSS.t1750 a_23564_n11428 a_21772_n11428.t1 VSS.t1749 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2173 VDD.t1583 a_46556_n12212 a_46468_n12168 VDD.t1582 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2174 a_33984_n10112 a_31872_n10529 a_33672_n10112 VDD.t3749 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X2175 a_13623_n14874.t2 a_21772_n11428.t13 VSS.t318 VSS.t317 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2176 VSS.t2911 a_33900_n11428 a_33364_n11384 VSS.t2910 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2177 a_2167_3472.t2 a_13623_n4162.t25 VSS.t580 VSS.t579 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2178 VSS.t2503 a_31279_n11728 a_31215_n11684 VSS.t2502 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2179 a_32359_n4372 a_33120_n3884 a_32911_n4240 VSS.t3642 nfet_06v0 ad=0.2007p pd=1.475u as=94.5f ps=0.885u w=0.36u l=0.6u
X2180 a_13501_n11816.t5 a_11023_n12196.t29 a_11087_n12816.t15 VDD.t131 pfet_03v3 ad=1.82p pd=6.9u as=0.728p ps=3.32u w=2.8u l=0.28u
X2181 VDD.t1811 a_37372_n10644 a_37284_n10600 VDD.t1810 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2182 VDD.t3723 a_28940_n2406.t5 a_30599_n12167 VDD.t3722 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2183 a_13501_n14494.t4 a_13623_n14874.t30 a_11087_n15494.t4 VSS.t1360 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2184 a_30451_n452 a_30781_n452 a_30901_n408 VSS.t3401 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X2185 a_13501_n17172.t14 a_11023_n17552.t30 a_11087_n18172.t14 VDD.t405 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2186 VSS.t2681 a_21692_n13308.t22 a_26532_n14437 VSS.t2680 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2187 a_37368_n320 a_35568_n4 a_36428_n53 VSS.t4091 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2188 a_23207_n4708 a_23887_n5156 VDD.t926 VDD.t925 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2189 a_30871_n11728 a_33910_n12146 VSS.t3622 VSS.t3621 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X2190 a_46668_n7941 a_46580_n7844 VSS.t3424 VSS.t3423 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2191 VDD.t1669 a_23564_n11428 a_21772_n11428.t6 VDD.t1668 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2192 a_24828_n18484 a_24740_n18440 VSS.t1669 VSS.t1668 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2193 VSS.t4013 a_30372_376 a_31076_376 VSS.t4012 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2194 a_43980_n4805 a_43892_n4708 VSS.t1986 VSS.t1985 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2195 a_26266_n9240 a_25642_n9816 a_26118_n9816 VSS.t2309 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2196 VDD.t1240 a_22588_n18917 a_22500_n18820 VDD.t1239 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2197 OUT[3].t7 a_38256_1564.t9 VSS.t174 VSS.t173 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2198 a_24041_816 a_24481_761.t50 a_24385_864 VSS.t796 nfet_06v0 ad=0.1989p pd=1.465u as=86.399994f ps=0.84u w=0.36u l=0.6u
X2199 a_36120_n4 a_35156_n325 a_35916_n4 VSS.t3065 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2200 a_23542_n1754 a_23954_n2020 a_24094_n1400 VDD.t2198 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2201 VDD.t3623 a_34649_n2412 a_25836_n1236.t6 VDD.t3622 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2202 VSS.t2691 a_26328_n6654.t18 a_21692_n13308.t1 VSS.t2690 nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2203 a_13501_n17172.t5 a_13623_n17552.t29 a_11087_n18172.t5 VSS.t88 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
D64 VSS.t513 a_23072_n13432.t60 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2204 a_37036_n9509 a_36948_n9412 VSS.t2356 VSS.t2355 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2205 VSS.t3157 a_33686_n11592 a_34162_n11593 VSS.t3156 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X2206 a_27744_n12908 a_21692_n13308.t23 VDD.t2621 VDD.t2620 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2207 a_37372_n16916 a_37284_n16872 VSS.t2939 VSS.t2938 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2208 VDD.t4267 a_46556_n5940 a_46468_n5896 VDD.t4266 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2209 a_27736_1248 a_25524_1243 a_26796_1515 VDD.t1365 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X2210 a_36252_n16916 a_36164_n16872 VSS.t3242 VSS.t3241 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2211 VDD.t512 a_23072_n13432.t61 a_30555_n13780 VDD.t511 pfet_06v0 ad=0.29465p pd=1.74u as=0.26p ps=1.52u w=1u l=0.5u
X2212 VDD.t983 a_46556_n2804 a_46468_n2760 VDD.t982 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2213 VSS.t798 a_24481_761.t51 a_42624_1248 VSS.t797 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2214 a_34392_n9815 a_25972_n6276 VSS.t1876 VSS.t1875 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X2215 a_11087_n15494.t30 a_2167_3472.t13 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X2216 VSS.t756 a_29800_n5940.t12 a_28156_n6412.t6 VSS.t755 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2217 a_34012_n16916 a_33924_n16872 VSS.t3182 VSS.t3181 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2218 a_43980_n15781 a_43892_n15684 VSS.t1919 VSS.t1918 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2219 a_22876_n1148 a_22568_n1104 VSS.t3009 VSS.t3008 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X2220 VDD.t1121 a_22876_n10556 a_22772_n10512 VDD.t1120 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2221 a_13501_n11816.t14 a_13623_n12196.t30 a_11087_n12816.t24 VSS.t1836 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2222 a_24578_n2020 a_24315_n2759 VSS.t3007 VSS.t3006 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2223 a_22876_n10556 a_22568_n10512 VDD.t1094 VDD.t1093 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X2224 a_41740_n15781 a_41652_n15684 VSS.t3084 VSS.t3083 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2225 a_13623_n4162.t1 a_21772_1116.t12 VSS.t473 VSS.t472 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2226 a_46556_n9076 a_46468_n9032 VSS.t4280 VSS.t4279 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2227 a_46108_n18484 a_46020_n18440 VSS.t3101 VSS.t3100 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2228 a_n263_3472.t10 a_22444_2253.t19 VDD.t2342 VDD.t457 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2229 a_44540_332 a_44452_376 VSS.t3284 VSS.t3283 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2230 a_40620_n15781 a_40532_n15684 VSS.t3234 VSS.t3233 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2231 VDD.t2496 a_44004_n1192 a_44640_1944.t4 VDD.t2495 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2232 a_22352_n12097 a_21940_n11684 VDD.t2190 VDD.t2189 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2233 a_46108_n15348 a_46020_n15304 VSS.t3068 VSS.t3067 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2234 a_43196_n13780 a_43108_n13736 VSS.t3624 VSS.t3623 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2235 VDD.t3912 a_43420_n1669 a_43332_n1572 VDD.t3911 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2236 a_29920_n12168 a_26388_n17606.t7 VDD.t237 VDD.t236 pfet_06v0 ad=0.224p pd=1.36u as=0.389p ps=2.02u w=0.56u l=0.5u
X2237 a_32650_n12168 a_32026_n12168 a_32482_n12168 VDD.t3705 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2238 a_43196_n10644 a_43108_n10600 VSS.t2333 VSS.t2332 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2239 a_43725_908 a_40260_n408 VDD.t2169 VDD.t2168 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X2240 VDD.t4287 a_47004_n15348 a_46916_n15304 VDD.t4286 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2241 a_45212_n2804 a_45124_n2760 VSS.t4352 VSS.t3293 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2242 VDD.t4291 a_48012_n6373 a_47924_n6276 VDD.t4290 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2243 VDD.t4293 a_37932_n15781 a_37844_n15684 VDD.t4292 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2244 VDD.t4295 a_48012_n3237 a_47924_n3140 VDD.t4294 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2245 a_11087_n23528.t19 a_11023_n22908.t30 a_13501_n22528.t15 VDD.t210 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2246 VDD.t3332 a_22876_n4284 a_22772_n4240 VDD.t3331 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2247 a_47564_n11077 a_47476_n10980 VSS.t1760 VSS.t1759 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2248 VDD.t4219 a_40060_n15348 a_39972_n15304 VDD.t4218 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2249 VSS.t2518 a_35849_n1192 a_36192_1248 VSS.t2517 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2250 a_26271_n1400 a_25647_n1976 a_26103_n1400 VDD.t1927 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2251 VSS.t3915 a_24771_n2804 a_24403_n2414 VSS.t3914 nfet_06v0 ad=0.14985p pd=1.145u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2252 a_31628_n5940.t8 a_33496_n6659.t20 VSS.t156 VSS.t155 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X2253 a_42636_n6373 a_42548_n6276 VSS.t2507 VSS.t2506 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2254 VDD.t3458 a_36812_n12645 a_36724_n12548 VDD.t3457 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2255 a_23024_n13248 a_22876_n13692 a_22856_n13248 VSS.t3928 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2256 VDD.t2206 a_26172_n20052 a_26084_n20008 VDD.t2205 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2257 VDD.t3707 a_47676_n20485 a_47588_n20388 VDD.t3706 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2258 a_35371_951 a_34895_376 a_35119_398 VSS.t2177 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X2259 a_24128_n704 a_21604_n708 a_23816_n704 VSS.t3435 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2260 a_34000_n3140 a_33588_n3461 VSS.t3422 VSS.t3421 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2261 a_21692_n5468.t5 a_26440_n5940.t10 VSS.t361 VSS.t360 nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X2262 VDD.t834 a_33776_n5896.t15 a_34708_n5896.t12 VDD.t833 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2263 a_42168_1564 a_41204_1243 a_41964_1564 VSS.t1870 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2264 a_45324_n11077 a_45236_n10980 VSS.t1201 VSS.t1200 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2265 VDD.t3492 a_45436_n20485 a_45348_n20388 VDD.t3491 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D65 VSS.t799 a_24481_761.t52 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2266 a_33496_n6659.t4 CLK.t7 VDD.t1821 VDD.t1820 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X2267 VSS.t4185 a_25940_n17606.t11 a_26299_n16388 VSS.t4184 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2268 a_38828_n15781 a_38740_n15684 VSS.t1022 VSS.t1021 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2269 a_22444_2253.t1 a_24236_2258.t7 VSS.t2441 VSS.t2440 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2270 a_23036_n16916 a_22948_n16872 VSS.t3788 VSS.t1871 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2271 VDD.t1608 a_24380_n18484 a_24292_n18440 VDD.t1607 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2272 VDD.t1080 a_25836_n1236.t16 a_29076_n8292.t0 VDD.t1079 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2273 OUT[1].t4 a_33216_1944.t16 VSS.t443 VSS.t442 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2274 VDD.t2690 a_24403_n2414 a_24315_n2759 VDD.t2689 pfet_06v0 ad=0.5346p pd=3.31u as=0.6561p ps=3.51u w=1.215u l=0.5u
X2275 VSS.t115 a_28156_n6412.t22 a_26328_n6654.t1 VSS.t114 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2276 VDD.t1610 a_22140_n18484 a_22052_n18440 VDD.t1609 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2277 a_24233_n8684 a_23072_n13432.t62 VDD.t514 VDD.t513 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X2278 a_11023_n17552.t15 a_13623_n17552.t30 VDD.t96 VDD.t95 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2279 a_28940_n2406.t0 a_29920_n3900.t16 a_31669_860 VSS.t654 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2280 VSS.t3773 a_28132_376 a_28836_376 VSS.t3772 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2281 a_27706_n1572 a_25836_n1236.t17 a_21916_n1975 VDD.t1081 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2282 VDD.t2463 a_38268_n15348 a_38180_n15304 VDD.t2462 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2283 a_38847_464 a_37947_332 VSS.t3370 VSS.t3369 nfet_06v0 ad=94.5f pd=0.885u as=0.1224p ps=1.04u w=0.36u l=0.6u
X2284 a_22568_n4240 a_22016_n4257 a_22364_n4240 VDD.t3265 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2285 VSS.t3544 a_37221_n3543 a_40196_n1884 VSS.t3543 nfet_06v0 ad=0.2344p pd=1.56u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2286 a_22892_n5156.t1 a_25237_n4327 a_32340_n5112 VSS.t1207 nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2287 a_37484_n9509 a_37396_n9412 VSS.t2877 VSS.t2876 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2288 a_22772_n10512 a_21604_n10116 a_22568_n10512 VDD.t3366 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2289 a_31961_n11340 a_31544_n11296 a_32337_n11296 VSS.t3124 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X2290 VDD.t3592 a_47900_n12212 a_47812_n12168 VDD.t3591 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2291 a_40280_864 a_39352_464 a_40112_864 VSS.t3301 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2292 a_39544_420 a_39056_820 a_39804_464 VDD.t948 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2293 VDD.t292 a_33496_n8222.t15 a_31548_n10172.t12 VDD.t291 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2294 a_11023_n12196.t10 a_13623_n12196.t31 VDD.t1750 VDD.t1749 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2295 a_41404_n9076 a_41316_n9032 VSS.t4146 VSS.t4145 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2296 a_11087_n23528.t43 a_2167_3472.t59 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X2297 a_27093_n7694 a_26973_n8292 VDD.t981 VDD.t980 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X2298 VDD.t1752 a_13623_n12196.t32 a_11023_n12196.t11 VDD.t1751 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2299 VSS.t758 a_29800_n5940.t13 a_28156_n6412.t5 VSS.t757 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2300 a_24760_n11383 a_25020_n11383 VSS.t1335 VSS.t1334 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X2301 a_36588_n11077 a_36500_n10980 VSS.t976 VSS.t975 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2302 VSS.t515 a_23072_n13432.t63 a_27952_n14432 VSS.t514 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2303 a_28076_n18484 a_27988_n18440 VSS.t1490 VSS.t1489 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2304 a_27820_n16432 a_24964_n14116 a_29479_n13735 VDD.t1837 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2305 VDD.t3391 a_25019_n3588.t5 a_29076_n8292.t3 VDD.t3390 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2306 a_11023_n14874.t10 a_13623_n14874.t31 VDD.t1310 VDD.t1309 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2307 VDD.t146 a_31628_n5940.t37 a_33776_n5896.t6 VDD.t145 pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X2308 a_27535_n12493 a_26635_n12996 VSS.t2128 VSS.t2127 nfet_06v0 ad=94.5f pd=0.885u as=0.1224p ps=1.04u w=0.36u l=0.6u
X2309 a_26499_n2732 a_25547_n2445 a_26935_n2272 VSS.t3976 nfet_06v0 ad=93.59999f pd=0.88u as=62.1f ps=0.705u w=0.36u l=0.6u
X2310 a_35800_n3456 a_33588_n3461 a_34860_n3189 VDD.t3338 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X2311 VDD.t3555 a_23932_n18917 a_23844_n18820 VDD.t3554 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2312 a_26944_n14116 a_26532_n14437 VDD.t1961 VDD.t1960 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2313 VSS.t582 a_13623_n4162.t26 a_2167_3472.t3 VSS.t581 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2314 VDD.t1452 a_37820_n5940 a_37732_n5896 VDD.t1451 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2315 a_13501_n9138.t3 a_11023_n9518.t27 a_11087_n10138.t7 VDD.t544 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2316 a_46220_n4805 a_46132_n4708 VSS.t2820 VSS.t2819 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2317 VDD.t3559 a_24604_n17349 a_24516_n17252 VDD.t3558 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D66 a_24481_761.t53 VDD.t738 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2318 a_44629_168 a_44509_n452 a_43885_n452 VDD.t1269 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2319 VSS.t403 a_21692_n5468.t22 a_21604_n708 VSS.t402 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2320 a_45660_n1236 a_45572_n1192 VSS.t2113 VSS.t2112 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2321 a_30616_n6221 a_30215_n6265 a_29559_n6456 VSS.t1887 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2322 VSS.t2521 a_26531_n10207 a_26239_n11428 VSS.t2520 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2323 a_39556_n4 a_38996_n408 a_39428_n408 VSS.t2488 nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X2324 VDD.t3926 a_25600_n5895 a_28583_n3140 VDD.t3925 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2325 a_36324_n4 a_35156_n325 a_36120_n4 VDD.t2986 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2326 VDD.t8 a_22444_332.t21 a_33252_n1192 VDD.t7 pfet_06v0 ad=0.4941p pd=2.03u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2327 a_45660_n2804 a_45572_n2760 VSS.t1560 VSS.t1559 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2328 a_35692_n18917 a_35604_n18820 VSS.t1301 VSS.t1300 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2329 VSS.t1093 a_21916_n6694.t10 a_28756_n5112 VSS.t1092 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2330 VDD.t1627 a_47900_n7508 a_47812_n7464 VDD.t1626 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2331 VDD.t2160 a_47116_n15781 a_47028_n15684 VDD.t2159 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2332 VDD.t2344 a_22444_2253.t20 a_n263_3472.t9 VDD.t2343 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2333 VDD.t1393 a_32262_n452 a_25940_n17606.t1 VDD.t1392 pfet_06v0 ad=0.4941p pd=2.03u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2334 a_41068_n5940 a_40980_n5896 VSS.t2987 VSS.t2986 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2335 VDD.t1482 a_47116_n12645 a_47028_n12548 VDD.t1481 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2336 VDD.t3426 a_41292_n15781 a_41204_n15684 VDD.t3425 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2337 a_24088_n16087 a_24348_n16087.t6 VSS.t2514 VSS.t1306 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X2338 VDD.t2224 a_29900_760.t10 a_38996_n408 VDD.t2223 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2339 a_23024_n704 a_22876_n1148 a_22856_n704 VSS.t2954 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2340 VDD.t2152 a_47900_n4372 a_47812_n4328 VDD.t2151 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2341 VDD.t330 a_10712_4516.t40 a_10778_2852.t6 VDD.t329 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2342 a_41292_n1669 a_41204_n1572 VSS.t4211 VSS.t4210 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2343 a_37820_n9076 a_37732_n9032 VSS.t2645 VSS.t2644 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2344 VDD.t2093 a_41292_n12645 a_41204_n12548 VDD.t2092 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2345 a_33452_n18917 a_33364_n18820 VSS.t2505 VSS.t2504 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2346 VDD.t1991 a_40172_n15781 a_40084_n15684 VDD.t1990 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2347 a_46220_n101 a_46132_n4 VSS.t972 VSS.t971 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2348 a_32332_n18917 a_32244_n18820 VSS.t1420 VSS.t1419 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2349 a_11087_n10138.t8 a_11023_n9518.t28 VSS.t561 VSS.t56 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2350 a_45660_n13780 a_45572_n13736 VSS.t3751 VSS.t3750 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2351 a_11087_n20850.t35 a_2167_3472.t22 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X2352 VSS.t1170 a_25084_1564 a_33216_1944.t0 VSS.t1169 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2353 a_31548_n10172.t11 a_33496_n8222.t16 VDD.t294 VDD.t293 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2354 a_45660_n10644 a_45572_n10600 VSS.t3354 VSS.t3353 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2355 VDD.t1985 a_35804_n12212 a_35716_n12168 VDD.t1984 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2356 a_44540_n13780 a_44452_n13736 VSS.t2203 VSS.t2202 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2357 VSS.t158 a_33496_n6659.t21 a_31628_n5940.t7 VSS.t157 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X2358 a_43555_n452 a_43885_n452 a_44005_n408 VSS.t4220 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X2359 a_33496_n6659.t5 CLK.t8 VDD.t1823 VDD.t1822 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X2360 a_44540_n10644 a_44452_n10600 VSS.t3161 VSS.t3160 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2361 a_23682_n1976 a_23542_n1754 a_22918_n2020 VSS.t2031 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X2362 a_29980_n5112 a_21916_n6694.t11 VSS.t1095 VSS.t1094 nfet_06v0 ad=0.1517p pd=1.19u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2363 a_21872_n12530 a_21996_n12996.t9 a_21892_n12952 VSS.t3575 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2364 a_42300_n13780 a_42212_n13736 VSS.t3534 VSS.t3533 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2365 VDD.t1464 a_30604_n11029 a_30500_n10980 VDD.t1463 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2366 a_42188_n15781 a_42100_n15684 VSS.t1406 VSS.t1405 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2367 a_43532_n9509 a_43444_n9412 VSS.t3238 VSS.t3237 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2368 a_42300_n10644 a_42212_n10600 VSS.t3303 VSS.t3302 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2369 a_26383_1944 a_25759_1944 a_26235_2520 VSS.t949 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2370 VDD.t2185 a_24716_1208.t2 a_24628_1252 VDD.t2184 pfet_06v0 ad=0.35315p pd=1.96u as=0.2486p ps=2.01u w=0.565u l=0.5u
X2371 a_39612_n4805 a_39524_n4708 VSS.t2568 VSS.t2567 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2372 a_34092_n9076 a_29532_n10311 VSS.t4064 VSS.t4063 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X2373 VDD.t4273 a_40956_n16916 a_40868_n16872 VDD.t4272 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2374 a_26328_n6654.t5 a_28156_n6412.t23 VDD.t124 VDD.t123 pfet_06v0 ad=0.2952p pd=1.54u as=0.367p ps=1.92u w=0.82u l=0.5u
X2375 VDD.t2143 a_25500_n10644 a_25412_n10600 VDD.t2142 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2376 VDD.t2527 a_40956_n13780 a_40868_n13736 VDD.t2526 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2377 a_11023_n6840.t9 a_13623_n6840.t30 VDD.t674 VDD.t673 pfet_03v3 ad=0.728p pd=3.32u as=1.82p ps=6.9u w=2.8u l=0.28u
X2378 a_34380_n408 a_29900_760.t11 a_34068_n4 VSS.t2298 nfet_06v0 ad=98.399994f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2379 a_28444_860 a_22444_332.t22 a_28132_376 VSS.t8 nfet_06v0 ad=98.399994f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2380 a_38256_1564.t2 a_37844_1564 VSS.t4264 VSS.t4263 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2381 VDD.t2107 a_41292_n6373 a_41204_n6276 VDD.t2106 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2382 a_35351_398 a_34895_376 a_35119_398 VDD.t2103 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X2383 VSS.t2551 a_40776_770 a_40672_864 VSS.t2550 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2384 VSS.t2339 a_28300_n15348 a_28849_n13252 VSS.t2338 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2385 VDD.t942 a_41292_n3237 a_41204_n3140 VDD.t941 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2386 a_40060_n4372 a_39972_n4328 VSS.t1241 VSS.t1240 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2387 a_40956_n20052 a_40868_n20008 VSS.t2228 VSS.t2227 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2388 VDD.t4130 a_32108_n2332.t22 a_35156_n325 VDD.t4129 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2389 VSS.t302 a_33496_n8222.t17 a_31548_n10172.t2 VSS.t301 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2390 a_41852_n9076 a_41764_n9032 VSS.t3226 VSS.t3225 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2391 VDD.t2623 a_21692_n13308.t24 a_22948_n14820 VDD.t2622 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2392 a_36155_n8548 a_25831_n11428 a_26172_n14564.t1 VSS.t1858 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2393 VDD.t887 a_23564_n20836 a_21772_n20836.t6 VDD.t886 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2394 a_38716_n18484 a_38628_n18440 VSS.t1635 VSS.t1634 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2395 a_29572_n5112 a_25836_n1236.t18 a_28548_n5112 VSS.t1108 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2396 VDD.t1639 a_29744_n15604.t16 a_23072_n13432.t5 VDD.t1638 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2397 VDD.t2625 a_21692_n13308.t25 a_26532_n14437 VDD.t2624 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2398 a_30452_n5156.t1 a_36744_n1954 VSS.t2875 VSS.t2874 nfet_06v0 ad=0.1261p pd=1.005u as=0.2134p ps=1.85u w=0.485u l=0.6u
X2399 a_27666_n5112 a_27190_n5112 a_27414_n5112 VSS.t1204 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X2400 a_38716_n15348 a_38628_n15304 VSS.t3078 VSS.t3077 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2401 a_34895_n1192 a_34271_n1192 a_34747_n616 VSS.t1402 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2402 VDD.t3934 a_30372_376 a_31076_376 VDD.t3933 pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X2403 a_47900_n1669 a_47812_n1572 VSS.t2717 VSS.t2716 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2404 a_31772_n18484 a_31684_n18440 VSS.t2555 VSS.t2554 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2405 VDD.t2651 a_47197_908 a_47317_376 VDD.t2650 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2406 a_24233_n3980 a_23816_n3840 a_24609_n3840 VSS.t2087 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X2407 VDD.t126 a_28156_n6412.t24 a_26328_n6654.t4 VDD.t125 pfet_06v0 ad=0.3608p pd=2.52u as=0.2952p ps=1.54u w=0.82u l=0.5u
X2408 VSS.t735 a_13623_n6840.t31 a_11023_n6840.t10 VSS.t734 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2409 VSS.t627 a_13623_n20230.t29 a_11023_n20230.t5 VSS.t626 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X2410 VSS.t3405 a_27452_n2716 a_27348_n2672 VSS.t3404 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2411 VSS.t1110 a_25836_n1236.t19 a_27628_n3841 VSS.t1109 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X2412 a_11023_n20230.t4 a_13623_n20230.t30 VSS.t629 VSS.t628 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2413 a_31856_1248 a_29332_1243 a_31544_1248 VSS.t2588 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2414 a_25559_n10980 a_26239_n11428 VDD.t964 VDD.t963 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2415 VDD.t3655 a_39612_n15348 a_39524_n15304 VDD.t3654 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2416 a_23228_n6679 a_21804_n2273.t7 a_23207_n4708 VDD.t1266 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2417 a_38156_n7941 a_38068_n7844 VSS.t2705 VSS.t2704 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D67 VSS.t835 a_22220_690.t10 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2418 VSS.t215 a_13623_n22908.t20 a_11023_n22908.t5 VSS.t214 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2419 a_31628_n5940.t26 a_33496_n6659.t22 VDD.t168 VDD.t167 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2420 a_11023_n22908.t4 a_13623_n22908.t21 VSS.t217 VSS.t216 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X2421 a_4001_4292.t0 a_3935_4156.t8 VSS.t458 VSS.t457 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X2422 a_38853_n1170 a_38733_n727 VDD.t1952 VDD.t1951 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X2423 a_39164_n7508 a_39076_n7464 VSS.t3209 VSS.t3208 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2424 VDD.t1198 a_33048_n7420 a_32856_n7376 VDD.t1197 pfet_06v0 ad=0.2222p pd=1.89u as=0.2424p ps=1.465u w=0.505u l=0.5u
X2425 a_13623_n17552.t12 a_21772_n8292.t16 VDD.t70 VDD.t69 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2426 a_4001_4292.t1 a_3935_4156.t9 a_3025_2852 VDD.t436 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X2427 VDD.t248 a_44640_1944.t14 OUT[5].t11 VDD.t247 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2428 VSS.t2269 a_24716_1208.t3 a_24628_1252 VSS.t2268 nfet_06v0 ad=0.2344p pd=1.56u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2429 VDD.t2531 a_29123_n6679 a_30900_n9032 VDD.t2530 pfet_06v0 ad=0.4941p pd=2.03u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2430 a_37932_n11077 a_37844_n10980 VSS.t4094 VSS.t4093 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2431 a_22788_n4708 a_21996_n12996.t10 a_22544_n4690 VDD.t3488 pfet_06v0 ad=0.3172p pd=1.74u as=0.4248p ps=1.94u w=1.22u l=0.5u
X2432 VDD.t3922 a_35064_1506 a_34872_1619 VDD.t3921 pfet_06v0 ad=0.2222p pd=1.89u as=0.2424p ps=1.465u w=0.505u l=0.5u
X2433 a_13501_n9138.t15 a_13623_n9518.t22 a_11087_n10138.t22 VSS.t253 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2434 VDD.t2047 a_36924_n20485 a_36836_n20388 VDD.t2046 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2435 VSS.t415 a_11023_n17552.t31 a_11087_n18172.t24 VSS.t68 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2436 VDD.t740 a_24481_761.t54 a_37947_332 VDD.t739 pfet_06v0 ad=0.29465p pd=1.74u as=0.26p ps=1.52u w=1u l=0.5u
X2437 VDD.t1444 a_44428_n7941 a_44340_n7844 VDD.t1443 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D68 VSS.t4137 a_22140_n6694.t10 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2438 VDD.t1989 a_26060_n18917 a_25972_n18820 VDD.t1988 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2439 a_38312_n1975 a_22276_n1572.t2 VDD.t4166 VDD.t4165 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X2440 a_29164_n5112 a_21916_n6694.t12 VSS.t1097 VSS.t1096 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2441 a_24573_n6724 a_22544_n4690 VDD.t2020 VDD.t2019 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X2442 a_11087_n10138.t21 a_13623_n9518.t23 a_13501_n9138.t14 VSS.t254 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X2443 VDD.t1139 a_46108_n12212 a_46020_n12168 VDD.t1138 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2444 VDD.t1003 a_35804_n20485 a_35716_n20388 VDD.t1002 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2445 a_28420_n14820 a_28300_n15348 VSS.t2337 VSS.t2336 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2446 VDD.t1501 a_44428_n4805 a_44340_n4708 VDD.t1500 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2447 a_30500_n10980 a_29332_n11301 a_30296_n10980 VDD.t3474 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2448 a_11087_n23528.t44 a_2167_3472.t58 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X2449 OUT[2].t6 a_37024_1944.t16 VSS.t1779 VSS.t1778 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2450 a_35288_n1975 a_32308_n1976 VDD.t3607 VDD.t3606 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X2451 VSS.t2523 a_38312_n1975 a_32636_n2020 VSS.t2522 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X2452 VDD.t2627 a_21692_n13308.t26 a_22052_n6980 VDD.t2626 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2453 a_26235_n3544 a_25759_n3544 VSS.t3569 VSS.t3568 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2454 a_30036_n7464 a_28736_n4633.t22 a_29888_n7464 VDD.t1035 pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X2455 a_33604_n5112 a_25836_n1236.t20 VSS.t1112 VSS.t1111 nfet_06v0 ad=0.1148p pd=1.1u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2456 VDD.t2102 a_39164_n10644 a_39076_n10600 VDD.t2101 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2457 VSS.t2714 a_32189_n9860 a_32309_n9816 VSS.t2713 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2458 a_23324_n7420 a_23016_n7376 VDD.t1494 VDD.t1493 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X2459 a_26643_n8292 a_26973_n8292 a_27093_n7694 VDD.t979 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2460 a_43980_n9509 a_43892_n9412 VSS.t2737 VSS.t2736 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2461 a_11087_n20850.t36 a_2167_3472.t23 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X2462 a_n263_3472.t1 a_22444_2253.t21 VSS.t2435 VSS.t2434 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2463 a_22672_n2759 a_21916_n1975 VDD.t1110 VDD.t1109 pfet_06v0 ad=0.44955p pd=1.955u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2464 VDD.t2028 a_47004_n9076 a_46916_n9032 VDD.t2027 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2465 VDD.t1736 a_27485_n10068 a_27605_n10600 VDD.t1735 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2466 a_25559_n12548 a_25831_n12996 a_25132_n16432 VDD.t2543 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2467 a_23404_816 a_25612_n878.t5 a_25524_n708 VSS.t846 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2468 a_22968_n6679 a_23228_n6679 VDD.t3243 VDD.t3242 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X2469 OUT[1].t3 a_33216_1944.t17 VSS.t445 VSS.t444 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2470 a_42188_n7941 a_42100_n7844 VSS.t3602 VSS.t3601 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2471 a_39164_n16916 a_39076_n16872 VSS.t3074 VSS.t3073 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2472 VSS.t882 a_33776_n5896.t16 a_34708_n5896.t2 VSS.t881 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2473 a_31628_n5940.t6 a_33496_n6659.t23 VSS.t160 VSS.t159 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X2474 a_2167_3472.t33 a_11023_n4162.t28 VSS.t2758 VDD.t2693 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2475 a_45324_n6373 a_45236_n6276 VSS.t2487 VSS.t2486 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D69 VSS.t4186 a_25940_n17606.t12 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2476 VSS.t3517 a_28153_1204 a_28048_1248 VSS.t3516 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X2477 VDD.t3430 a_26060_n878.t2 a_23404_816 VDD.t3429 pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X2478 a_13623_n20230.t4 a_21772_n3588.t12 VSS.t912 VSS.t911 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2479 VDD.t4215 a_21692_n15348 a_21604_n15304 VDD.t1787 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2480 a_32413_n14564 a_28752_n15348 VSS.t3203 VSS.t3202 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2481 a_27452_n2716 a_28736_1944 a_28791_n3543 VSS.t1280 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2482 a_43196_n7508 a_43108_n7464 VSS.t3940 VSS.t3939 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2483 a_45772_n15781 a_45684_n15684 VSS.t4152 VSS.t4151 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2484 VDD.t3284 a_37947_332 a_37859_377 VDD.t3283 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2485 a_34428_n452.t0 a_37785_n364 VSS.t1903 VSS.t1902 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2486 VDD.t1436 a_42076_n2804 a_41988_n2760 VDD.t1435 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2487 a_13501_n14494.t14 a_11023_n14874.t30 a_11087_n15494.t14 VDD.t78 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2488 a_27884_332.t0 a_29519_n1976 VSS.t2417 VSS.t2416 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X2489 a_39357_n660 a_30732_332.t3 VSS.t1687 VSS.t1686 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2490 VSS.t2300 a_29900_760.t12 a_41684_n1976 VSS.t2299 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2491 a_28617_n8548 a_28721_n9076.t7 a_28225_n9031 VDD.t415 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2492 VSS.t3072 a_28232_n12606 a_28040_n12493 VSS.t3071 nfet_06v0 ad=0.2016p pd=1.48u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2493 a_13623_n9518.t3 a_21772_n17700.t12 VDD.t1009 VDD.t1008 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2494 a_43532_n15781 a_43444_n15684 VSS.t4177 VSS.t4176 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2495 a_28548_n5112 a_24815_n3588.t14 a_31788_n5112 VSS.t23 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2496 a_13623_n12196.t13 a_21772_n14564.t8 VDD.t2006 VDD.t2005 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2497 a_33815_1384 a_34576_1204 a_34367_1619 VSS.t1641 nfet_06v0 ad=0.2007p pd=1.475u as=94.5f ps=0.885u w=0.36u l=0.6u
X2498 VDD.t3816 a_23703_n5156.t2 a_25559_n10980 VDD.t3815 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2499 a_43196_n18484 a_43108_n18440 VSS.t1639 VSS.t1638 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2500 a_31455_n13648 a_30555_n13780 VSS.t1712 VSS.t1711 nfet_06v0 ad=94.5f pd=0.885u as=0.1224p ps=1.04u w=0.36u l=0.6u
X2501 a_24264_n6976 a_22052_n6980 a_23324_n7420 VDD.t1489 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X2502 VDD.t3998 a_25948_n20485 a_25860_n20388 VDD.t3997 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2503 VSS.t3222 a_25817_804 a_25769_860 VSS.t3221 nfet_06v0 ad=0.14985p pd=1.145u as=48.6f ps=0.645u w=0.405u l=0.6u
X2504 a_28972_n8247 a_28852_n8292.t2 a_28764_n8247 VSS.t3667 nfet_06v0 ad=0.2119p pd=1.335u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2505 a_13501_n17172.t13 a_11023_n17552.t32 a_11087_n18172.t13 VDD.t406 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2506 a_43196_n15348 a_43108_n15304 VSS.t3917 VSS.t3916 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2507 VDD.t3697 a_28132_376 a_28836_376 VDD.t3696 pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X2508 VDD.t3635 a_39724_n9509 a_39636_n9412 VDD.t3634 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2509 VSS.t3431 a_25627_n452 a_25539_n407.t0 VSS.t3430 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2510 a_38403_n5503 a_38733_n5431 a_38853_n5321 VSS.t2243 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X2511 a_45212_n7508 a_45124_n7464 VSS.t2001 VSS.t2000 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2512 VSS.t1526 a_26736_n364 a_26631_7 VSS.t1525 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2513 a_28009_n12168 a_27279_n12146 VSS.t2614 VSS.t2613 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X2514 a_34142_n12146 a_33686_n11592 a_33910_n12146 VDD.t3076 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X2515 VDD.t1633 a_44092_n15348 a_44004_n15304 VDD.t1632 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2516 VSS.t134 a_31628_n5940.t38 a_29800_n5940.t0 VSS.t133 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2517 VDD.t2043 a_39724_n15781 a_39636_n15684 VDD.t2042 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2518 a_25817_804 a_24913_864 VSS.t3011 VSS.t3010 nfet_06v0 ad=0.1782p pd=1.69u as=0.14985p ps=1.145u w=0.405u l=0.6u
X2519 a_22016_n1121 a_21604_n708 VDD.t3359 VDD.t3358 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2520 a_36388_n1572 a_35940_n1931 VDD.t3027 VDD.t3026 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
D70 VSS.t516 a_23072_n13432.t64 diode_nd2ps_06v0 pj=1.86u area=0.2052p
D71 VSS.t1309 a_21804_n2273.t8 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2521 a_13501_n11816.t4 a_11023_n12196.t30 a_11087_n12816.t14 VDD.t132 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2522 a_11087_n15494.t5 a_13623_n14874.t32 a_13501_n14494.t5 VSS.t1361 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2523 a_31628_n5940.t25 a_33496_n6659.t24 VDD.t170 VDD.t169 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
D72 a_22140_n6694.t11 VDD.t4063 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2524 OUT[4].t8 a_41392_1944.t15 VDD.t1387 VDD.t1386 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2525 VDD.t3605 a_31961_1204 a_31856_1248 VDD.t3604 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X2526 VSS.t2759 a_11023_n4162.t29 VSS.t2759 VSS.t64 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.28u
X2527 VDD.t2085 a_38604_n12645 a_38516_n12548 VDD.t2084 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2528 VSS.t2145 a_26383_1944 a_26859_2519 VSS.t2144 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X2529 a_10778_2852.t6 a_10712_4516.t41 VDD.t332 VDD.t331 pfet_03v3 ad=0.728p pd=3.32u as=1.82p ps=6.9u w=2.8u l=0.28u
X2530 VSS.t3137 a_40196_1944 a_41392_1944.t3 VSS.t3136 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2531 VSS.t518 a_23072_n13432.t65 a_23024_n3840 VSS.t517 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2532 VDD.t676 a_13623_n6840.t32 a_11023_n6840.t11 VDD.t675 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2533 VDD.t10 a_22444_332.t23 a_33900_n11428 VDD.t9 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X2534 a_47116_n11077 a_47028_n10980 VSS.t2804 VSS.t2803 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2535 VDD.t2738 a_27988_n20388 a_30192_n15304.t5 VDD.t2737 pfet_06v0 ad=0.367p pd=1.92u as=0.2952p ps=1.54u w=0.82u l=0.5u
X2536 VDD.t2096 a_25573_n12167 a_28225_n9031 VDD.t415 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2537 VDD.t1458 a_47228_n20485 a_47140_n20388 VDD.t1457 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2538 a_41292_n11077 a_41204_n10980 VSS.t3765 VSS.t3764 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D73 VSS.t800 a_24481_761.t55 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2539 VDD.t968 a_44876_n7941 a_44788_n7844 VDD.t967 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2540 a_26527_51 a_25627_n452 VSS.t3429 VSS.t3428 nfet_06v0 ad=94.5f pd=0.885u as=0.1224p ps=1.04u w=0.36u l=0.6u
X2541 a_39477_n1192 a_39357_n660 a_38733_n727 VDD.t2133 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2542 a_40172_n11077 a_40084_n10980 VSS.t2834 VSS.t2833 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2543 VDD.t894 a_44876_n4805 a_44788_n4708 VDD.t893 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2544 VDD.t2113 a_37372_n7508 a_37284_n7464 VDD.t2112 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2545 a_31909_n12952 a_31789_n12996 VSS.t4360 VSS.t4359 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X2546 a_34796_n15781 a_34708_n15684 VSS.t1915 VSS.t1914 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2547 VSS.t644 a_21772_1116.t13 a_13623_n4162.t0 VSS.t643 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2548 a_11087_n7460.t16 a_11023_n6840.t30 VSS.t107 VSS.t58 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2549 VDD.t1143 a_26172_n18484 a_26084_n18440 VDD.t1142 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2550 VDD.t2350 a_24236_2258.t8 a_22444_2253.t4 VDD.t2349 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2551 a_11087_n12816.t25 a_13623_n12196.t33 a_13501_n11816.t15 VSS.t1837 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2552 OUT[5].t10 a_44640_1944.t15 VDD.t250 VDD.t249 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2553 a_28144_n4708 a_27414_n5112 VSS.t3919 VSS.t3918 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X2554 VDD.t558 a_13623_n4162.t27 a_11023_n4162.t16 VDD.t557 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2555 VDD.t742 a_24481_761.t56 a_25627_n452 VDD.t741 pfet_06v0 ad=0.29465p pd=1.74u as=0.26p ps=1.52u w=1u l=0.5u
X2556 VDD.t2120 a_47452_n9076 a_47364_n9032 VDD.t2119 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2557 a_46220_n18917 a_46132_n18820 VSS.t3148 VSS.t3147 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2558 a_47004_n1236 a_46916_n1192 VSS.t4325 VSS.t4324 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2559 VSS.t584 a_13623_n4162.t28 a_2167_3472.t4 VSS.t583 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2560 VDD.t3231 a_24731_n3124.t3 a_26060_n878.t0 VDD.t3230 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X2561 a_45772_n6373 a_45684_n6276 VSS.t2529 VSS.t2528 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2562 VSS.t2437 a_22444_2253.t22 a_n263_3472.t0 VSS.t2436 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
D74 a_22220_690.t11 VDD.t782 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2563 a_10778_2852.t3 a_10712_4516.t42 VDD.t334 VDD.t333 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2564 a_39648_n2020 a_26553_377.t4 VSS.t129 VSS.t128 nfet_06v0 ad=0.1584p pd=1.6u as=0.2344p ps=1.56u w=0.36u l=0.6u
X2565 VDD.t1041 a_30452_n5156.t6 a_28736_n4633.t12 VDD.t1040 pfet_06v0 ad=0.4056p pd=1.805u as=0.2197p ps=1.365u w=0.845u l=0.5u
D75 a_24481_761.t57 VDD.t743 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2566 VSS.t1221 a_23564_n8292 a_21772_n8292.t2 VSS.t1220 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2567 VDD.t2156 a_40956_n20052 a_40868_n20008 VDD.t2155 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2568 a_22140_n15781 a_22052_n15684 VSS.t4214 VSS.t4126 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2569 a_29199_n3543 a_25600_n5895 a_27452_n2716 VSS.t4007 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X2570 a_46220_n9509 a_46132_n9412 VSS.t1545 VSS.t1544 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2571 a_22096_376 a_22220_690.t12 a_22116_860 VSS.t472 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2572 VSS.t1689 a_30732_332.t4 a_30684_860 VSS.t1688 nfet_06v0 ad=0.2132p pd=1.34u as=98.399994f ps=1.06u w=0.82u l=0.6u
X2573 a_39556_n4 a_29900_760.t13 a_39408_n4 VDD.t2225 pfet_06v0 ad=0.3172p pd=1.74u as=0.1464p ps=1.46u w=1.22u l=0.5u
X2574 VDD.t4190 a_37844_1564 a_38256_1564.t6 VDD.t4189 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2575 a_22876_n1148 a_22568_n1104 VDD.t2933 VDD.t2932 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X2576 a_33851_n1976 a_33375_n1976 VSS.t2028 VSS.t2027 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2577 a_45660_n7508 a_45572_n7464 VSS.t4021 VSS.t4020 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2578 a_11087_n20850.t37 a_2167_3472.t24 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X2579 VDD.t991 a_41516_n5940 a_41428_n5896 VDD.t990 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2580 a_31965_n8292 a_29123_n6679 VDD.t2529 VDD.t2528 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X2581 VDD.t3771 a_45212_332 a_45124_376 VDD.t3770 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2582 a_24264_n6976 a_22464_n7393 a_23324_n7420 VSS.t4115 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2583 a_28764_n8247 a_29076_n8292.t8 a_28972_n8247 VSS.t469 nfet_06v0 ad=0.4137p pd=1.9u as=0.2119p ps=1.335u w=0.815u l=0.6u
X2584 a_33900_n11428 a_30871_n11728 VDD.t896 VDD.t895 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X2585 a_37484_n18917 a_37396_n18820 VSS.t1874 VSS.t1873 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2586 a_26266_n13736 a_25642_n13736 a_26098_n13736 VDD.t1183 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2587 a_21772_n3588.t2 a_23564_n3588.t5 VSS.t2993 VSS.t2992 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2588 VSS.t1192 a_39357_n5364 a_39477_n5320 VSS.t1191 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2589 a_36520_n3868 a_10712_4516.t43 VDD.t336 VDD.t335 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X2590 a_29900_n10600.t0 a_29444_n10116 VSS.t2039 VSS.t2038 nfet_06v0 ad=0.3608p pd=2.52u as=0.2344p ps=1.56u w=0.82u l=0.6u
D76 VSS.t9 a_22444_332.t24 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2591 VDD.t1983 a_43084_n15781 a_42996_n15684 VDD.t1982 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2592 a_42556_n1976 a_29900_760.t14 a_42244_n1572 VSS.t2301 nfet_06v0 ad=98.399994f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2593 a_41180_n2804 a_41092_n2760 VSS.t982 VSS.t981 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2594 VSS.t520 a_23072_n13432.t66 a_30752_n11296 VSS.t519 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2595 a_24693_n12376 a_24573_n12996 a_23949_n12996 VDD.t2587 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2596 VDD.t1424 a_43084_n12645 a_42996_n12548 VDD.t1423 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2597 a_35244_n18917 a_35156_n18820 VSS.t3861 VSS.t3860 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2598 a_28492_n12548 a_28040_n12493 VDD.t3773 VDD.t3772 pfet_06v0 ad=0.2028p pd=1.3u as=0.45p ps=2.02u w=0.78u l=0.5u
X2599 a_27852_n14990 a_28121_n10980 VDD.t3599 VDD.t3598 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X2600 a_44540_n9076 a_44452_n9032 VSS.t2419 VSS.t2418 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2601 a_45660_n18484 a_45572_n18440 VSS.t3950 VSS.t3949 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2602 VDD.t3188 a_38716_n12212 a_38628_n12168 VDD.t3187 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2603 a_44540_n18484 a_44452_n18440 VSS.t2907 VSS.t2906 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2604 a_45660_n15348 a_45572_n15304 VSS.t2871 VSS.t2870 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2605 a_47452_n13780 a_47364_n13736 VSS.t1516 VSS.t1515 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2606 a_39428_n408 a_39308_n452 VSS.t2733 VSS.t2732 nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2607 VSS.t866 a_34708_n5896.t23 a_33496_n8222.t1 VSS.t865 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2608 VSS.t2760 a_11023_n4162.t30 a_2167_3472.t34 VDD.t2694 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2609 a_47452_n10644 a_47364_n10600 VSS.t2883 VSS.t2882 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2610 a_44540_n15348 a_44452_n15304 VSS.t3325 VSS.t3324 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2611 a_32132_n4708 a_25237_n4327 a_22892_n5156.t0 VDD.t1168 pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2612 VDD.t1967 a_30320_n6636 a_30215_n6265 VDD.t1966 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2613 a_29056_n14432 a_26532_n14437 a_28744_n14432 VSS.t2035 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2614 VDD.t1942 a_37859_377 a_39760_n4 VDD.t1941 pfet_06v0 ad=0.4392p pd=1.94u as=0.4758p ps=2u w=1.22u l=0.5u
X2615 a_42300_n18484 a_42212_n18440 VSS.t1988 VSS.t1987 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2616 a_45212_n13780 a_45124_n13736 VSS.t1652 VSS.t1651 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2617 VDD.t1854 a_34068_n4 a_34403_332 VDD.t1853 pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X2618 a_35568_n4 a_35156_n325 VSS.t3064 VSS.t3063 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2619 a_42300_n15348 a_42212_n15304 VSS.t3412 VSS.t3411 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2620 a_44428_n3237 a_44340_n3140 VSS.t3396 VSS.t3395 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2621 VDD.t2360 a_42300_n9076 a_42212_n9032 VDD.t2359 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2622 a_45212_n10644 a_45124_n10600 VSS.t3224 VSS.t3223 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2623 a_28153_1204 a_24481_761.t58 VDD.t745 VDD.t744 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X2624 VDD.t2298 a_42748_n16916 a_42660_n16872 VDD.t2297 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2625 VDD.t2162 a_42771_769 a_40776_770 VDD.t2161 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2626 VDD.t1862 a_24233_n3980 a_24128_n3840 VDD.t1861 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X2627 VDD.t2409 a_23999_n2320.t5 a_25647_n1976 VDD.t2408 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2628 VDD.t2722 a_42748_n13780 a_42660_n13736 VDD.t2721 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D77 a_24481_761.t59 VDD.t746 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2629 a_29180_n9387 a_26388_n17606.t8 a_28868_n9387 VDD.t238 pfet_06v0 ad=0.2847p pd=1.615u as=0.58035p ps=2.155u w=1.095u l=0.5u
X2630 VDD.t2653 a_40508_n16916 a_40420_n16872 VDD.t2652 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2631 a_42771_769 a_43101_841 a_43221_398 VDD.t1850 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2632 a_22568_n4240 a_21604_n3844 a_22364_n4240 VSS.t1805 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2633 VSS.t522 a_23072_n13432.t67 a_27123_n12872 VSS.t521 nfet_06v0 ad=0.1224p pd=1.04u as=0.134p ps=1.1u w=0.36u l=0.6u
X2634 VDD.t1680 a_40508_n13780 a_40420_n13736 VDD.t1679 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2635 a_32351_n7376 a_31451_n7508 VSS.t4248 VSS.t4247 nfet_06v0 ad=94.5f pd=0.885u as=0.1224p ps=1.04u w=0.36u l=0.6u
X2636 VDD.t4206 a_22220_n12996 a_22116_n12548 VDD.t4205 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2637 a_21772_1116.t2 a_23564_1116.t6 VSS.t3497 VSS.t3496 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2638 VSS.t4246 a_31451_n7508 a_25020_n8200.t0 VSS.t4245 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2639 a_30807_n11684 a_27988_n4328 VSS.t1577 VSS.t1576 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2640 a_29856_n1121 a_29444_n708 VDD.t2744 VDD.t2743 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2641 VDD.t252 a_44640_1944.t16 OUT[5].t9 VDD.t251 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2642 a_11087_n10138.t9 a_11023_n9518.t29 VSS.t562 VSS.t58 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2643 a_42748_n20052 a_42660_n20008 VSS.t2392 VSS.t2391 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2644 a_29751_n1422 a_29295_n1400 a_29519_n1976 VDD.t1485 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X2645 VDD.t1893 a_24672_n11339 a_24836_n4708 VDD.t1892 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2646 VDD.t2381 a_47116_n7941 a_47028_n7844 VDD.t2380 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2647 a_29744_1564 a_29332_1243 VSS.t2587 VSS.t2586 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2648 a_26727_n1422 a_26271_n1400 a_26495_n1976 VDD.t2507 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X2649 VDD.t2392 a_47116_n4805 a_47028_n4708 VDD.t2391 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2650 VSS.t4167 a_35456_n4628.t16 a_32108_n2332.t2 VSS.t4166 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2651 a_40508_n20052 a_40420_n20008 VSS.t2380 VSS.t2379 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2652 VSS.t2153 a_32152_n13692 a_31960_n13648 VSS.t2152 nfet_06v0 ad=0.2016p pd=1.48u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2653 VDD.t947 a_39056_820 a_38951_420 VDD.t946 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2654 a_35392_n10172 a_34652_n11391 VDD.t4153 VDD.t4152 pfet_06v0 ad=0.2486p pd=2.01u as=0.35315p ps=1.96u w=0.565u l=0.5u
X2655 VDD.t3702 XRST.t2 a_27540_n20747 VDD.t3701 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X2656 VDD.t2148 a_35692_n13780 a_35604_n13736 VDD.t2147 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2657 a_32308_n1572 a_29532_n4372.t5 VDD.t2053 VDD.t2052 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2658 a_33900_n15781 a_33812_n15684 VSS.t2479 VSS.t2478 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2659 OUT[1].t2 a_33216_1944.t18 VSS.t447 VSS.t446 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2660 a_42096_n1572 a_37859_377 VDD.t1940 VDD.t1939 pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2661 VSS.t3139 a_30036_n7464 a_30740_n7464 VSS.t3138 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2662 a_29540_n11728 a_29532_n10311 VSS.t4062 VSS.t4061 nfet_06v0 ad=0.176p pd=1.68u as=0.104p ps=0.92u w=0.4u l=0.6u
X2663 VDD.t3330 a_33488_n12996 a_23564_n14564.t1 VDD.t3329 pfet_06v0 ad=0.35315p pd=1.96u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2664 VDD.t397 a_21692_n5468.t23 a_25524_1243 VDD.t396 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2665 a_33564_n18484 a_33476_n18440 VSS.t1152 VSS.t1151 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2666 a_27195_n6889 a_26719_n7464 a_26943_n7442 VSS.t2532 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X2667 a_25831_n11428 a_27526_n9816 VDD.t2375 VDD.t2374 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X2668 a_33077_n1191 a_32073_n844 VSS.t3099 VSS.t3098 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2669 a_11023_n14874.t11 a_13623_n14874.t33 VSS.t1363 VSS.t1362 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2670 a_35849_n1192 a_35119_n1170 VSS.t2925 VSS.t2924 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X2671 a_43420_n1669 a_43332_n1572 VSS.t3994 VSS.t3856 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2672 a_31324_n18484 a_31236_n18440 VSS.t2164 VSS.t2163 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2673 a_26571_n6888 a_26095_n7464 VSS.t1161 VSS.t1160 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2674 a_21692_2431 a_28153_1204 VSS.t3515 VSS.t3514 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2675 VSS.t1114 a_25836_n1236.t21 a_31676_n3544 VSS.t1113 nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X2676 a_42372_1564 a_41204_1243 a_42168_1564 VDD.t1783 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2677 VDD.t2702 a_41964_n5940 a_41876_n5896 VDD.t2701 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2678 VSS.t90 a_13623_n17552.t31 a_11023_n17552.t4 VSS.t89 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X2679 a_22672_n2759 a_23004_n2332 a_22672_n2214.t1 VDD.t3590 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2680 a_33416_n4240 a_33120_n3884 a_32359_n4372 VDD.t3553 pfet_06v0 ad=0.2424p pd=1.465u as=0.25375p ps=1.51u w=0.505u l=0.5u
X2681 a_48012_n6373 a_47924_n6276 VSS.t4354 VSS.t4353 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2682 a_11023_n17552.t3 a_13623_n17552.t32 VSS.t92 VSS.t91 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2683 a_36324_n4 a_24481_761.t60 VDD.t748 VDD.t747 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X2684 a_44004_n1192 a_43556_n661 VSS.t1384 VSS.t1383 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X2685 a_39724_n11077 a_39636_n10980 VSS.t3460 VSS.t3459 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2686 a_22856_n704 a_22016_n1121 a_22568_n1104 VSS.t3439 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2687 VDD.t1929 a_30716_n1148 a_30612_n1104 VDD.t1928 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2688 VSS.t176 a_38256_1564.t10 OUT[3].t6 VSS.t175 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2689 a_43555_n452 a_43885_n452 a_44005_146 VDD.t4147 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2690 a_29652_n3844 a_29532_n4372.t6 VSS.t2123 VSS.t2122 nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2691 VDD.t4098 a_38716_n20485 a_38628_n20388 VDD.t2192 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2692 VSS.t1740 a_36388_1944 a_37024_1944.t2 VSS.t1739 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2693 a_11087_n10138.t10 a_11023_n9518.t30 a_13501_n9138.t4 VDD.t545 pfet_03v3 ad=0.728p pd=3.32u as=1.82p ps=6.9u w=2.8u l=0.28u
X2694 VSS.t868 a_34708_n5896.t24 a_33496_n8222.t0 VSS.t867 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2695 a_32502_n11592 a_32026_n12168 VSS.t3778 VSS.t3777 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2696 VDD.t1213 a_43196_n12212 a_43108_n12168 VDD.t1212 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2697 a_11023_n12196.t12 a_13623_n12196.t34 VSS.t1839 VSS.t1838 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2698 VDD.t612 a_29920_n3900.t17 a_24815_n3588.t2 VDD.t611 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2699 VDD.t4119 a_25940_n17606.t13 a_25412_n5895 VDD.t4118 pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X2700 a_25972_n6276 a_25524_n6635 VSS.t3382 VSS.t3381 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X2701 VDD.t1522 a_30652_n20485 a_30564_n20388 VDD.t1521 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2702 VDD.t2883 a_35848_n3868 a_23564_n3588.t1 VDD.t2882 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2703 a_44876_n12645 a_44788_n12548 VSS.t3844 VSS.t3843 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2704 a_44876_n3237 a_44788_n3140 VSS.t3180 VSS.t3179 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2705 a_24698_n1400 a_24578_n2020 a_23954_n2020 VDD.t4224 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2706 VDD.t3195 a_24681_n7116 a_24576_n6976 VDD.t3194 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X2707 a_13623_n14874.t15 a_21772_n11428.t14 VDD.t302 VDD.t301 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2708 a_42636_n12645 a_42548_n12548 VSS.t1609 VSS.t1608 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2709 VSS.t3135 a_40196_1944 a_41392_1944.t2 VSS.t3134 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2710 a_31936_n6592 a_30320_n6636 a_30808_n6334 VSS.t2047 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2711 a_23038_n1976 a_22918_n2020 VSS.t4111 VSS.t4110 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X2712 VDD.t3508 a_30584_n1954 a_21996_n12996.t2 VDD.t3507 pfet_06v0 ad=0.458p pd=2.02u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2713 VDD.t2475 a_35392_n10172 a_28519_n10160.t1 VDD.t2474 pfet_06v0 ad=0.35315p pd=1.96u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2714 a_22588_n18484 a_22500_n18440 VSS.t3787 VSS.t3786 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2715 VSS.t3374 a_39556_n4 a_40260_n408 VSS.t3373 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2716 a_23016_n7376 a_22052_n6980 a_22812_n7376 VSS.t1553 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
D78 VSS.t10 a_22444_332.t25 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2717 a_28156_n6412.t11 a_29800_n5940.t14 VDD.t700 VDD.t699 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2718 a_30408_n1104 a_29856_n1121 a_30204_n1104 VDD.t944 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2719 a_22444_332.t3 a_27259_804.t11 VDD.t803 VDD.t802 pfet_06v0 ad=0.52205p pd=2.045u as=0.4334p ps=2.85u w=0.985u l=0.5u
X2720 VSS.t2308 a_24684_n16432 a_22600_n12124 VSS.t2307 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X2721 VDD.t4002 a_28300_n20485 a_28212_n20388 VDD.t4001 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2722 a_24348_n16087.t1 a_25577_n14956 VDD.t2826 VDD.t2825 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2723 a_47564_n15781 a_47476_n15684 VSS.t2289 VSS.t2288 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2724 VSS.t3759 a_30900_n9032 a_21692_n6694.t0 VSS.t3758 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2725 OUT[5].t8 a_44640_1944.t17 VDD.t274 VDD.t273 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2726 a_24771_n2804 a_25795_n2716.t3 a_25139_n2704 VSS.t2451 nfet_06v0 ad=93.59999f pd=0.88u as=0.2898p ps=2.33u w=0.36u l=0.6u
X2727 VDD.t2292 a_47564_n7941 a_47476_n7844 VDD.t2291 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2728 VSS.t219 a_13623_n22908.t22 a_11023_n22908.t3 VSS.t218 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2729 a_21772_n17700.t6 a_23564_n17700 VDD.t4247 VDD.t4246 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2730 a_36192_1248 a_34576_1204 a_35064_1506 VSS.t1640 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2731 VDD.t2183 a_47564_n4805 a_47476_n4708 VDD.t2182 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2732 VDD.t2394 a_36364_n7941 a_36276_n7844 VDD.t2393 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2733 a_45324_n15781 a_45236_n15684 VSS.t2773 VSS.t2772 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2734 a_47452_n1236 a_47364_n1192 VSS.t2413 VSS.t2412 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2735 VSS.t4169 a_35456_n4628.t17 a_32108_n2332.t1 VSS.t4168 nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2736 VDD.t1011 a_21772_n17700.t13 a_13623_n9518.t4 VDD.t1010 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2737 a_21772_n14564.t1 a_23564_n14564.t4 VDD.t3740 VDD.t3739 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2738 VSS.t4293 a_24578_n2020 a_24698_n1976 VSS.t4292 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2739 a_29732_n2760 a_27259_804.t12 a_27628_n3841 VDD.t804 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2740 VDD.t1919 a_21772_n14564.t9 a_13623_n12196.t12 VDD.t1918 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2741 VSS.t1781 a_37024_1944.t17 OUT[2].t5 VSS.t1780 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2742 a_22968_n6679 a_23228_n6679 VSS.t3329 VSS.t3328 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X2743 VDD.t2256 a_44876_n17349 a_44788_n17252 VDD.t2255 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2744 a_40112_864 a_24481_761.t61 VSS.t802 VSS.t801 nfet_06v0 ad=43.199997f pd=0.6u as=0.2016p ps=1.48u w=0.36u l=0.6u
X2745 a_47317_952 a_47197_908 a_46573_841 VSS.t2708 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X2746 a_30111_n6221 a_29211_n6724 VDD.t3960 VDD.t3959 pfet_06v0 ad=0.1313p pd=1.025u as=0.29465p ps=1.74u w=0.505u l=0.5u
X2747 VDD.t2316 a_44876_n14213 a_44788_n14116 VDD.t2315 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2748 a_31968_n704 a_29444_n708 a_31656_n704 VSS.t2817 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2749 VDD.t930 a_39648_n2020 a_23564_1116.t1 VDD.t929 pfet_06v0 ad=0.35315p pd=1.96u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2750 a_22016_n8961 a_21604_n8548 VDD.t3953 VDD.t3952 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
D79 VSS.t836 a_22220_690.t13 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2751 VDD.t2373 a_42636_n17349 a_42548_n17252 VDD.t2372 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2752 a_48012_n101 a_47924_n4 VSS.t2313 VSS.t2312 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2753 a_22016_n5825 a_21604_n5412 VDD.t3495 VDD.t3494 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2754 a_21812_n6276 a_21692_n6694.t19 VDD.t640 VDD.t364 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2755 VDD.t1083 a_25836_n1236.t22 a_24631_n3588 VDD.t1082 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2756 a_27597_n8292 a_24716_n5156.t5 VDD.t1327 VDD.t1326 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X2757 a_11087_n20850.t24 a_13623_n20230.t31 a_13501_n19850.t14 VSS.t630 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2758 VSS.t2443 a_24236_2258.t9 a_22444_2253.t0 VSS.t2442 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2759 a_11087_n7460.t15 a_11023_n6840.t31 VSS.t108 VSS.t66 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2760 a_24604_n17349 a_24516_n17252 VSS.t948 VSS.t947 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2761 VDD.t2643 a_42636_n14213 a_42548_n14116 VDD.t2642 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2762 a_24965_n9860 a_25724_n14564 a_25636_n14520 VSS.t3042 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2763 VDD.t2367 a_35692_n15781 a_35604_n15684 VDD.t2366 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2764 VSS.t449 a_33216_1944.t19 OUT[1].t1 VSS.t448 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2765 a_27852_n18917 a_27764_n18820 VSS.t3211 VSS.t3210 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2766 a_10778_2852.t4 a_10712_4516.t44 VSS.t349 VSS.t348 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2767 a_34727_n1192 a_34271_n1192 VDD.t1348 VDD.t1347 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X2768 VDD.t2296 a_34572_n12645 a_34484_n12548 VDD.t2295 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2769 a_11087_n23528.t5 a_13623_n22908.t23 a_13501_n22528.t5 VSS.t220 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2770 VDD.t3992 a_33452_n15781 a_33364_n15684 VDD.t3144 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2771 a_30604_1515 a_30296_1564 VSS.t3654 VSS.t3653 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X2772 a_30472_n9815 a_28617_n8548 VDD.t2596 VDD.t2595 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X2773 a_25612_n18917 a_25524_n18820 VSS.t2181 VSS.t2180 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2774 a_11023_n6840.t12 a_13623_n6840.t33 VSS.t737 VSS.t736 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2775 a_31548_n10172.t10 a_33496_n8222.t18 VDD.t296 VDD.t295 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2776 a_39477_n5896 a_39357_n5364 a_38733_n5431 VDD.t1146 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2777 a_43084_n11077 a_42996_n10980 VSS.t4029 VSS.t4028 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2778 a_25831_n12996 a_27526_n13714 VSS.t2306 VSS.t2305 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X2779 a_29540_n11728 a_29532_n10311 a_30180_n12168 VDD.t3982 pfet_06v0 ad=0.2464p pd=2u as=0.1736p ps=1.18u w=0.56u l=0.5u
X2780 VDD.t2245 a_26755_n16132 a_26239_n12996 VDD.t2244 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2781 a_39477_n2760 a_39357_n2228 a_38733_n2295 VDD.t2763 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2782 a_34756_n3140 a_24481_761.t62 VDD.t750 VDD.t749 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X2783 VDD.t2736 a_27988_n20388 a_30192_n15304.t4 VDD.t761 pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X2784 a_37820_n13780 a_37732_n13736 VSS.t1589 VSS.t1588 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2785 VSS.t3703 a_34649_n2412 a_25836_n1236.t0 VSS.t3702 nfet_06v0 ad=0.3586p pd=2.51u as=0.2119p ps=1.335u w=0.815u l=0.6u
X2786 a_37820_n10644 a_37732_n10600 VSS.t3305 VSS.t3304 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2787 VSS.t670 a_21772_n20836.t16 a_13623_n6840.t1 VSS.t669 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2788 VDD.t3979 a_42076_n20485 a_41988_n20388 VDD.t3978 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2789 a_28752_n15348 a_29161_n14476 VSS.t2745 VSS.t2744 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2790 a_27988_n20388 a_27540_n20747 VDD.t2878 VDD.t2877 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X2791 a_36588_n15781 a_36500_n15684 VSS.t1034 VSS.t1033 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2792 VDD.t2666 a_40396_n7941 a_40308_n7844 VDD.t2665 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2793 a_13623_n6840.t0 a_21772_n20836.t17 VSS.t672 VSS.t671 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2794 a_29900_760.t1 a_33252_n1192 VDD.t1275 VDD.t1274 pfet_06v0 ad=0.3782p pd=1.84u as=0.4941p ps=2.03u w=1.22u l=0.5u
X2795 VDD.t4021 a_44092_n7508 a_44004_n7464 VDD.t4020 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2796 VDD.t881 a_31011_n8292 a_30396_n7508 VDD.t880 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2797 a_11087_n15494.t31 a_2167_3472.t12 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X2798 a_34348_n15781 a_34260_n15684 VSS.t1773 VSS.t1772 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2799 a_11087_n15494.t13 a_11023_n14874.t31 a_13501_n14494.t13 VDD.t79 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2800 VDD.t3418 a_44092_n4372 a_44004_n4328 VDD.t3417 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2801 a_28968_n12864 a_28040_n12493 a_28800_n12864 VSS.t3849 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2802 VDD.t806 a_27259_804.t13 a_25612_n878.t0 VDD.t805 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X2803 VDD.t3970 a_44204_n5940 a_44116_n5896 VDD.t3969 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2804 a_31936_n6592 a_30215_n6265 a_30808_n6334 VDD.t1806 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2805 a_21872_n12530 a_21772_n12996 VDD.t3639 VDD.t3638 pfet_06v0 ad=0.4248p pd=1.94u as=0.4972p ps=3.14u w=1.13u l=0.5u
X2806 a_48012_n18917 a_47924_n18820 VSS.t2928 VSS.t2927 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2807 VSS.t524 a_23072_n13432.t68 a_31043_n13248 VSS.t523 nfet_06v0 ad=0.1224p pd=1.04u as=0.134p ps=1.1u w=0.36u l=0.6u
X2808 a_27167_n10808 a_26543_n11384 a_27019_n11384 VSS.t2020 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
D80 a_22140_n6694.t12 VDD.t4064 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2809 VDD.t1576 a_30988_n18917 a_30900_n18820 VDD.t1575 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2810 a_29263_n3588.t0 a_27225_n1572.t2 VDD.t3480 VDD.t3479 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X2811 VDD.t353 a_26440_n5940.t11 a_21692_n5468.t11 VDD.t352 pfet_06v0 ad=0.367p pd=1.92u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2812 VSS.t320 a_21772_n11428.t15 a_13623_n14874.t1 VSS.t319 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2813 VDD.t2925 a_24152_n11680 a_24569_n11820 VDD.t2924 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X2814 VDD.t2726 a_45660_n12212 a_45572_n12168 VDD.t2725 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2815 VDD.t3660 a_23564_n452.t3 a_21772_n452.t1 VDD.t3659 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2816 VDD.t264 a_13623_n9518.t24 a_11023_n9518.t14 VDD.t263 pfet_03v3 ad=1.82p pd=6.9u as=0.728p ps=3.32u w=2.8u l=0.28u
X2817 a_13623_n14874.t0 a_21772_n11428.t16 VSS.t322 VSS.t321 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2818 a_33126_n11592 a_32650_n12168 a_32854_n12168 VSS.t3269 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X2819 VDD.t3942 a_44540_n12212 a_44452_n12168 VDD.t3941 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2820 VDD.t1283 a_27672_n3543 a_21692_n7508.t1 VDD.t1282 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2821 a_41292_n6373 a_41204_n6276 VSS.t2117 VSS.t2116 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2822 a_23304_n6976 a_22464_n7393 a_23016_n7376 VSS.t4114 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2823 VDD.t338 a_10712_4516.t45 a_10778_2852.t7 VDD.t337 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2824 OUT[4].t7 a_41392_1944.t16 VSS.t1428 VSS.t1427 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2825 a_40672_864 a_38951_420 a_39544_420 VDD.t3217 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2826 VDD.t2263 a_42604_n2020 a_42448_n1572 VDD.t2262 pfet_06v0 ad=0.4392p pd=1.94u as=0.4758p ps=2u w=1.22u l=0.5u
X2827 VSS.t2321 a_23507_n2759 a_25423_n4328 VSS.t2320 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X2828 a_11087_n12816.t13 a_11023_n12196.t31 a_13501_n11816.t3 VDD.t133 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2829 a_26503_n4306 a_26047_n4328 a_26271_n4306 VDD.t2592 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X2830 a_26981_n10578 a_26861_n10135 VDD.t1542 VDD.t1541 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X2831 VDD.t1708 a_42300_n12212 a_42212_n12168 VDD.t1707 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2832 a_11023_n4162.t5 a_13623_n4162.t29 VSS.t586 VSS.t585 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2833 a_47116_n3237 a_47028_n3140 VSS.t3121 VSS.t3120 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2834 a_28156_n6412.t4 a_29800_n5940.t15 VSS.t760 VSS.t759 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2835 VDD.t2306 a_42748_n20052 a_42660_n20008 VDD.t2305 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2836 a_10712_4516.t24 a_10778_2852.t26 VDD.t377 VDD.t376 pfet_03v3 ad=0.728p pd=3.32u as=1.82p ps=6.9u w=2.8u l=0.28u
X2837 a_22876_n8988 a_22568_n8944 VDD.t3670 VDD.t3669 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X2838 a_26172_n14564.t0 a_25831_n11428 VDD.t1772 VDD.t1771 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X2839 VSS.t3879 a_42244_n1572 a_42948_n1976 VSS.t3878 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2840 a_37708_n7941 a_37620_n7844 VSS.t1284 VSS.t1283 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2841 VDD.t304 a_21772_n11428.t17 a_13623_n14874.t14 VDD.t303 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2842 a_23932_n18484 a_23844_n18440 VSS.t2224 VSS.t2223 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2843 VSS.t2761 a_11023_n4162.t31 a_2167_3472.t35 VDD.t2695 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2844 a_22876_n5852 a_22568_n5808 VDD.t1026 VDD.t1025 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X2845 a_31068_n6276 a_30616_n6221 VDD.t2122 VDD.t2121 pfet_06v0 ad=0.2028p pd=1.3u as=0.45p ps=2.02u w=0.78u l=0.5u
D81 a_21804_n2273.t9 VDD.t1267 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2846 VDD.t4016 a_40508_n20052 a_40420_n20008 VDD.t4015 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2847 VDD.t909 a_21692_n18917 a_21604_n18820 VDD.t908 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2848 VSS.t1047 a_21772_n17700.t14 a_13623_n9518.t5 VSS.t1046 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2849 VDD.t1825 a_47452_1900 a_47364_1944 VDD.t1824 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2850 a_24578_n2020 a_24315_n2759 VDD.t2931 VDD.t2930 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
D82 VSS.t4187 a_25940_n17606.t14 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2851 a_27829_n16088 a_27709_n16132 a_27085_n16132 VSS.t3589 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X2852 VSS.t1991 a_21772_n14564.t10 a_13623_n12196.t5 VSS.t1990 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2853 a_46693_398 a_46573_841 VDD.t2732 VDD.t2731 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X2854 a_33999_n1400 a_33375_n1976 a_33851_n1976 VSS.t2026 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2855 a_29559_n6456 a_30320_n6636 a_30111_n6221 VSS.t2046 nfet_06v0 ad=0.2007p pd=1.475u as=94.5f ps=0.885u w=0.36u l=0.6u
X2856 a_25472_n14816 a_22948_n14820 a_25160_n14816 VSS.t2108 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2857 a_38716_n7508 a_38628_n7464 VSS.t1211 VSS.t1210 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2858 a_39276_n18917 a_39188_n18820 VSS.t3207 VSS.t3206 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2859 VDD.t1141 a_25237_n13735 a_25642_n13736 VDD.t1140 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2860 VSS.t405 a_21692_n5468.t24 a_21604_n5412 VSS.t404 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2861 VDD.t3440 a_40956_n18484 a_40868_n18440 VDD.t3439 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2862 VDD.t225 a_13623_n22908.t24 a_11023_n22908.t15 VDD.t224 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2863 VDD.t3268 a_44316_n1236 a_44228_n1192 VDD.t3068 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2864 a_11023_n22908.t14 a_13623_n22908.t25 VDD.t227 VDD.t226 pfet_03v3 ad=0.728p pd=3.32u as=1.82p ps=6.9u w=2.8u l=0.28u
X2865 a_37036_n18917 a_36948_n18820 VSS.t3268 VSS.t3267 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2866 a_23642_n1400 a_23542_n1754 a_22918_n2020 VDD.t1958 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2867 a_26859_2519 a_26383_1944 a_26607_1966 VSS.t2143 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X2868 a_47452_n18484 a_47364_n18440 VSS.t3695 VSS.t3694 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2869 a_47004_n4372 a_46916_n4328 VSS.t3613 VSS.t3612 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2870 a_36388_1944 a_35940_2475 VSS.t3524 VSS.t3523 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X2871 a_30092_n18917 a_30004_n18820 VSS.t3256 VSS.t3255 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2872 a_47452_n15348 a_47364_n15304 VSS.t2721 VSS.t2720 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2873 a_45212_n18484 a_45124_n18440 VSS.t4322 VSS.t4321 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2874 VDD.t399 a_21692_n5468.t25 a_21604_n3844 VDD.t398 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2875 VSS.t687 a_21692_n6694.t20 a_34092_n9076 VSS.t686 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2876 a_40060_n9076 a_39972_n9032 VSS.t2626 VSS.t2625 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2877 VSS.t369 a_26440_n5940.t12 a_21692_n5468.t4 VSS.t368 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2878 a_45212_n15348 a_45124_n15304 VSS.t2725 VSS.t2724 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2879 a_47004_n13780 a_46916_n13736 VSS.t4006 VSS.t4005 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2880 VDD.t340 a_10712_4516.t46 a_10778_2852.t8 VDD.t339 pfet_03v3 ad=1.82p pd=6.9u as=0.728p ps=3.32u w=2.8u l=0.28u
X2881 a_47004_n10644 a_46916_n10600 VSS.t2933 VSS.t2932 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2882 a_11087_n20850.t38 a_2167_3472.t26 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X2883 VSS.t2762 a_11023_n4162.t32 VSS.t2762 VSS.t56 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.28u
X2884 VSS.t4189 a_25940_n17606.t15 a_36155_n8548 VSS.t4188 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2885 a_13501_n19850.t4 a_11023_n20230.t30 a_11087_n20850.t10 VDD.t1847 pfet_03v3 ad=1.82p pd=6.9u as=0.728p ps=3.32u w=2.8u l=0.28u
X2886 a_40060_n13780 a_39972_n13736 VSS.t4052 VSS.t4051 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2887 VDD.t1995 CLK.t9 a_33496_n6659.t4 VDD.t1994 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X2888 a_27605_n10024 a_27485_n10068 a_26861_n10135 VSS.t1815 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X2889 a_40060_n10644 a_39972_n10600 VSS.t3661 VSS.t3660 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D83 VSS.t803 a_24481_761.t63 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2890 a_23415_n5111 a_21804_n2273.t10 VSS.t1311 VSS.t1310 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2891 VSS.t1099 a_21916_n6694.t13 a_29572_n5112 VSS.t1098 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2892 VDD.t172 a_33496_n6659.t25 a_31628_n5940.t24 VDD.t171 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2893 a_44988_n20485 a_44900_n20388 VSS.t4119 VSS.t4118 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2894 a_43868_n20485 a_43780_n20388 VSS.t3292 VSS.t3291 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2895 VSS.t1738 a_36388_1944 a_37024_1944.t1 VSS.t1737 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2896 OUT[3].t14 a_38256_1564.t11 VDD.t192 VDD.t191 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2897 a_32108_n2332.t11 a_35456_n4628.t18 VDD.t4089 VDD.t4088 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2898 a_25732_n1192 a_25612_n878.t6 VDD.t797 VDD.t796 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X2899 VSS.t256 a_13623_n9518.t25 a_11023_n9518.t4 VSS.t255 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2900 VDD.t1562 a_46780_n20485 a_46692_n20388 VDD.t1561 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2901 a_26531_n10207 a_26861_n10135 a_26981_n10025 VSS.t1620 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X2902 VDD.t2089 a_32158_n12212 a_32026_n12168 VDD.t2088 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2903 VDD.t3414 a_43833_1204 a_43728_1248 VDD.t3413 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X2904 a_24233_n844 a_23072_n13432.t69 VDD.t516 VDD.t515 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X2905 a_42748_n7508 a_42660_n7464 VSS.t2409 VSS.t2408 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2906 a_27758_n9262 a_27302_n9816 a_27526_n9816 VDD.t1930 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X2907 a_41628_n20485 a_41540_n20388 VSS.t3803 VSS.t3802 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2908 VDD.t586 a_13623_n20230.t32 a_11023_n20230.t15 VDD.t585 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2909 VDD.t3304 a_41628_n2804 a_41540_n2760 VDD.t3303 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2910 a_22772_n10512 a_23072_n13432.t70 VDD.t518 VDD.t517 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X2911 a_28247_n10599 a_28927_n10160 VDD.t2312 VDD.t2311 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2912 VSS.t109 a_11023_n6840.t32 a_11087_n7460.t14 VSS.t68 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2913 VDD.t1294 a_44540_n20485 a_44452_n20388 VDD.t1293 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2914 a_11023_n20230.t14 a_13623_n20230.t33 VDD.t588 VDD.t587 pfet_03v3 ad=0.728p pd=3.32u as=1.82p ps=6.9u w=2.8u l=0.28u
X2915 VDD.t952 a_43420_n20485 a_43332_n20388 VDD.t951 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2916 VDD.t1085 a_25836_n1236.t23 a_29444_n4328.t2 VDD.t1084 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X2917 a_21812_n6643 a_22140_n6694.t13 VSS.t4138 VSS.t2672 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X2918 a_37932_n15781 a_37844_n15684 VSS.t4356 VSS.t4355 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2919 a_13623_n6840.t13 a_21772_n20836.t18 VDD.t624 VDD.t623 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2920 a_22140_n16916 a_22052_n16872 VSS.t4127 VSS.t4126 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2921 VDD.t2678 a_40508_n7508 a_40420_n7464 VDD.t2677 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2922 a_25139_n2704 a_24403_n2414 VDD.t2688 VDD.t2687 pfet_06v0 ad=0.2028p pd=1.3u as=0.3276p ps=1.62u w=0.78u l=0.5u
X2923 a_23816_n3840 a_21604_n3844 a_22876_n4284 VDD.t1715 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X2924 VDD.t1456 a_40508_n4372 a_40420_n4328 VDD.t1455 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2925 a_31011_n8292 a_31341_n8292 a_31461_n8248 VSS.t4048 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X2926 VDD.t2660 a_41740_n9509 a_41652_n9412 VDD.t2659 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2927 a_35356_n18484 a_35268_n18440 VSS.t1716 VSS.t1715 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2928 a_47564_n3237 a_47476_n3140 VSS.t3258 VSS.t3257 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2929 a_28156_n6412.t3 a_29800_n5940.t16 VSS.t762 VSS.t761 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2930 a_28121_n10980 a_27391_n11384 VSS.t3683 VSS.t3682 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X2931 VDD.t3258 a_35244_n13780 a_35156_n13736 VDD.t1368 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2932 a_38268_n13780 a_38180_n13736 VSS.t3553 VSS.t3552 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2933 a_28548_n5112 a_25836_n1236.t24 a_29164_n5112 VSS.t1115 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2934 a_38268_n10644 a_38180_n10600 VSS.t4068 VSS.t4067 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2935 VSS.t2583 a_26271_n1400 a_26747_n1976 VSS.t2582 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X2936 VDD.t3410 a_23564_1116.t7 a_21772_1116.t3 VDD.t2345 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2937 a_33116_n18484 a_33028_n18440 VSS.t4025 VSS.t4024 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2938 VSS.t3641 a_33120_n3884 a_33015_n4284 VSS.t3640 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2939 VDD.t752 a_24481_761.t64 a_33308_n7376 VDD.t751 pfet_06v0 ad=0.45p pd=2.02u as=0.3432p ps=2.44u w=0.78u l=0.5u
X2940 a_39724_n9509 a_39636_n9412 VSS.t3723 VSS.t3722 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2941 VDD.t1191 a_37372_n15348 a_37284_n15304 VDD.t1190 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2942 VSS.t1430 a_41392_1944.t17 OUT[4].t6 VSS.t1429 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2943 a_33955_1240 a_33815_1384 a_33467_1116 VSS.t1041 nfet_06v0 ad=0.134p pd=1.1u as=0.176p ps=1.68u w=0.4u l=0.6u
X2944 a_38853_n2185 a_38733_n2295 VSS.t2825 VSS.t2824 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X2945 VDD.t2116 a_27628_n18484 a_27540_n18440 VDD.t2115 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2946 a_27348_n2672 a_25795_n2716.t4 a_26499_n2732 VSS.t2452 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2947 a_24573_n12996 a_21872_n12530 VSS.t1945 VSS.t1944 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2948 a_11087_n20850.t39 a_2167_3472.t27 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X2949 a_35816_n174 a_35119_398 VDD.t419 VDD.t418 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X2950 a_42157_n660 a_34428_n452.t6 VSS.t3052 VSS.t3051 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2951 VSS.t1117 a_25836_n1236.t25 a_34372_n5112 VSS.t1116 nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
D84 a_24481_761.t65 VDD.t753 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2952 VSS.t351 a_10712_4516.t47 a_10778_2852.t9 VSS.t350 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2953 VDD.t3896 a_29408_1944.t16 OUT[0].t15 VDD.t3895 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2954 VDD.t755 a_24481_761.t66 a_35324_1564 VDD.t754 pfet_06v0 ad=0.45p pd=2.02u as=0.3432p ps=2.44u w=0.78u l=0.5u
X2955 a_37632_n2020 a_36388_n1572 VSS.t1069 VSS.t1068 nfet_06v0 ad=0.1584p pd=1.6u as=0.2344p ps=1.56u w=0.36u l=0.6u
X2956 VSS.t902 a_25020_n8200.t3 a_29532_n10311 VSS.t901 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X2957 VDD.t808 a_27259_804.t14 a_29444_n4328.t1 VDD.t807 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X2958 VSS.t2648 a_26047_n4328 a_26523_n3753 VSS.t2647 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X2959 a_27180_n18484 a_27092_n18440 VSS.t4009 VSS.t4008 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2960 a_47452_n4372 a_47364_n4328 VSS.t3820 VSS.t3819 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2961 a_13623_n17552.t2 a_21772_n8292.t17 VSS.t53 VSS.t52 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2962 VSS.t2115 a_30676_n7844 a_31919_n9032 VSS.t2114 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X2963 VDD.t4073 a_39052_n7941 a_38964_n7844 VDD.t4072 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2964 a_32581_n9860 a_28435_n10599 a_33364_n11384 VSS.t3168 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2965 VDD.t1163 a_33564_n20485 a_33476_n20388 VDD.t1162 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2966 a_34544_n2272 a_32432_n2689 a_34232_n2272 VDD.t3389 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X2967 a_27778_n9816 a_27302_n9816 a_27526_n9816 VSS.t3377 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X2968 a_26175_n11383 a_23703_n5156.t3 a_24684_n16432 VSS.t3897 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X2969 VDD.t2068 a_32444_n20485 a_32356_n20388 VDD.t2067 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2970 a_24069_n12952 a_23949_n12996 VSS.t1250 VSS.t1249 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X2971 a_46668_n12645 a_46580_n12548 VSS.t2867 VSS.t2866 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2972 a_27784_n14432 a_26944_n14116 a_27496_n14116 VSS.t3999 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2973 VDD.t757 a_24481_761.t67 a_27484_n4 VDD.t756 pfet_06v0 ad=0.45p pd=2.02u as=0.3432p ps=2.44u w=0.78u l=0.5u
X2974 VSS.t451 a_33216_1944.t20 OUT[1].t0 VSS.t450 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2975 a_32911_n4240 a_31787_n3969 VDD.t1528 VDD.t1527 pfet_06v0 ad=0.1313p pd=1.025u as=0.33755p ps=1.955u w=0.505u l=0.5u
X2976 a_24069_n6680 a_23949_n6724 VSS.t989 VSS.t988 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X2977 a_11023_n14874.t12 a_13623_n14874.t34 VSS.t1365 VSS.t1364 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2978 a_47900_n2804 a_47812_n2760 VSS.t2837 VSS.t2716 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2979 a_44428_n12645 a_44340_n12548 VSS.t1706 VSS.t1705 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2980 VSS.t1975 a_11023_n20230.t31 a_11087_n20850.t11 VSS.t70 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2981 VDD.t1170 a_30204_n20485 a_30116_n20388 VDD.t1169 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2982 a_32888_n13248 a_31960_n13648 a_32720_n13248 VSS.t3614 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2983 VSS.t2208 a_39357_n660 a_39477_n616 VSS.t2207 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2984 a_24752_n16132 a_24716_n5156.t6 VSS.t1378 VSS.t1377 nfet_06v0 ad=0.1584p pd=1.6u as=0.2344p ps=1.56u w=0.36u l=0.6u
X2985 a_35351_n1170 a_34895_n1192 a_35119_n1170 VDD.t1395 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X2986 a_40396_n3237 a_40308_n3140 VSS.t2979 VSS.t2978 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2987 a_43308_n5940 a_43220_n5896 VSS.t3639 VSS.t3638 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2988 a_30616_n6221 a_30320_n6636 a_29559_n6456 VDD.t1965 pfet_06v0 ad=0.2424p pd=1.465u as=0.25375p ps=1.51u w=0.505u l=0.5u
X2989 VDD.t2648 a_39500_n6373 a_39412_n6276 VDD.t2647 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2990 a_11087_n20850.t12 a_11023_n20230.t32 VSS.t1976 VSS.t72 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X2991 a_11087_n23528.t45 a_2167_3472.t57 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X2992 VDD.t1100 a_46220_n15781 a_46132_n15684 VDD.t1099 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2993 VSS.t178 a_38256_1564.t12 OUT[3].t5 VSS.t177 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2994 a_31324_n4372 a_31348_n1931 VDD.t1102 VDD.t1101 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X2995 VSS.t1905 a_23619_n6724 a_22264_n5852 VSS.t1904 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2996 VDD.t2563 a_28437_n13705 a_28247_n10599 VDD.t2562 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2997 VDD.t1161 a_39500_n3237 a_39412_n3140 VDD.t1160 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2998 VDD.t4202 a_46220_n12645 a_46132_n12548 VDD.t4201 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2999 a_32579_769 a_32909_841 a_33029_398 VDD.t4250 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
D85 a_23072_n13432.t71 VDD.t519 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3000 a_34089_n10252 a_33672_n10112 a_34465_n10112 VSS.t3549 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X3001 a_26887_n12168 a_26431_n12168 VDD.t3176 VDD.t3175 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X3002 a_21772_n9860 a_23479_n5156 VDD.t2239 VDD.t2238 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X3003 VDD.t278 a_31548_n10172.t21 a_31460_n10116 VDD.t277 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X3004 a_28756_n5112 a_25836_n1236.t26 a_28548_n5112 VSS.t1118 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3005 VSS.t162 a_33496_n6659.t26 a_31628_n5940.t5 VSS.t161 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X3006 a_39056_820 a_32108_n2332.t23 VDD.t4132 VDD.t4131 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X3007 a_11023_n12196.t13 a_13623_n12196.t35 VSS.t1841 VSS.t1840 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3008 a_47116_n15781 a_47028_n15684 VSS.t1756 VSS.t1755 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3009 OUT[2].t4 a_37024_1944.t18 VSS.t1783 VSS.t1782 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3010 a_40956_n12212 a_40868_n12168 VSS.t2956 VSS.t2955 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3011 a_11087_n23528.t23 a_11023_n22908.t31 VSS.t198 VSS.t56 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3012 VDD.t4245 a_23564_n17700 a_21772_n17700.t5 VDD.t4244 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3013 VDD.t4182 a_40956_n7508 a_40868_n7464 VDD.t4181 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3014 VDD.t4184 a_43084_n7941 a_42996_n7844 VDD.t4183 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3015 a_41292_n15781 a_41204_n15684 VSS.t3713 VSS.t3712 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3016 a_13623_n9518.t6 a_21772_n17700.t15 VDD.t1013 VDD.t1012 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3017 a_40172_n15781 a_40084_n15684 VSS.t2070 VSS.t2069 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3018 VDD.t3742 a_23564_n14564.t5 a_21772_n14564.t2 VDD.t3741 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3019 VDD.t3615 a_40956_n4372 a_40868_n4328 VDD.t3614 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3020 VDD.t3794 a_43084_n4805 a_42996_n4708 VDD.t3793 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3021 VDD.t3709 a_44876_n18917 a_44788_n18820 VDD.t3708 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3022 VDD.t4164 a_46668_n17349 a_46580_n17252 VDD.t4163 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3023 VDD.t1015 a_21772_n17700.t16 a_13623_n9518.t3 VDD.t1014 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3024 a_13623_n12196.t11 a_21772_n14564.t11 VDD.t1921 VDD.t1920 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3025 VDD.t4178 a_46668_n14213 a_46580_n14116 VDD.t4177 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3026 VDD.t1874 a_21772_n14564.t12 a_13623_n12196.t10 VDD.t1873 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3027 VSS.t3298 a_41336_n407 a_24236_2258.t0 VSS.t3297 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X3028 VSS.t2873 a_36744_n1954 a_30452_n5156.t0 VSS.t2872 nfet_06v0 ad=0.151p pd=1.185u as=0.1261p ps=1.005u w=0.485u l=0.6u
X3029 a_35025_n2272 a_24481_761.t68 VSS.t805 VSS.t804 nfet_06v0 ad=0.217p pd=1.515u as=0.1224p ps=1.04u w=0.36u l=0.6u
X3030 a_27175_n7442 a_26719_n7464 a_26943_n7442 VDD.t2454 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X3031 VDD.t1499 a_42636_n18917 a_42548_n18820 VDD.t1498 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3032 VDD.t4151 a_44428_n17349 a_44340_n17252 VDD.t4150 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3033 a_31909_n14520 a_31789_n14564 VSS.t2561 VSS.t2560 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X3034 a_13623_n20230.t10 a_21772_n3588.t13 VDD.t859 VDD.t858 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3035 VDD.t84 a_21772_n8292.t18 a_13623_n17552.t11 VDD.t83 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3036 a_10778_2852.t12 a_4001_4292.t9 VSS.t892 VSS.t354 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3037 a_36192_1248 a_34471_1575 a_35064_1506 VDD.t3957 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3038 VDD.t4168 a_44428_n14213 a_44340_n14116 VDD.t4167 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3039 VSS.t2030 a_23542_n1754 a_23682_n1976 VSS.t2029 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3040 a_40732_n2804 a_40644_n2760 VSS.t2800 VSS.t2799 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3041 VDD.t2447 a_43532_n6373 a_43444_n6276 VDD.t2446 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3042 VSS.t2917 a_27055_n12168 a_27531_n11593 VSS.t2916 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X3043 VDD.t4159 a_37484_n15781 a_37396_n15684 VDD.t4158 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3044 a_13501_n14494.t6 a_13623_n14874.t35 a_11087_n15494.t6 VSS.t1366 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3045 VDD.t2150 a_43532_n3237 a_43444_n3140 VDD.t2149 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3046 a_42300_n4372 a_42212_n4328 VSS.t2142 VSS.t2141 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3047 a_29644_n18917 a_29556_n18820 VSS.t3088 VSS.t3087 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3048 a_26944_1248 a_26796_1515 a_26776_1248 VSS.t2580 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3049 a_34756_n3140 a_33588_n3461 a_34552_n3140 VDD.t3337 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3050 VDD.t2062 a_36364_n12645 a_36276_n12548 VDD.t2061 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3051 VDD.t954 a_35244_n15781 a_35156_n15684 VDD.t953 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3052 OUT[1].t10 a_33216_1944.t21 VDD.t431 VDD.t430 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
D86 a_22444_332.t26 VDD.t11 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3053 a_11087_n18172.t4 a_13623_n17552.t33 a_13501_n17172.t4 VSS.t93 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3054 a_35848_n3868 a_25237_n4327 VDD.t1167 VDD.t1166 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X3055 a_24180_n5112 a_24492_n5156 VSS.t3586 VSS.t3585 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3056 VDD.t148 a_31628_n5940.t39 a_33776_n5896.t5 VDD.t147 pfet_06v0 ad=0.367p pd=1.92u as=0.2952p ps=1.54u w=0.82u l=0.5u
X3057 a_24233_n10252 a_23816_n10112 a_24609_n10112 VSS.t2007 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X3058 a_31760_n12168 a_30787_n12167 VSS.t1907 VSS.t1906 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X3059 a_27404_n18917 a_27316_n18820 VSS.t3753 VSS.t3752 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D87 a_24481_761.t69 VDD.t758 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3060 VSS.t3659 a_27167_n10808 a_27643_n11384 VSS.t3658 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X3061 VDD.t626 a_21772_n20836.t19 a_13623_n6840.t12 VDD.t625 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3062 a_37820_n18484 a_37732_n18440 VSS.t2160 VSS.t2159 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3063 a_38161_n320 a_24481_761.t70 VSS.t807 VSS.t806 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X3064 a_32911_n4240 a_31787_n3969 VSS.t1593 VSS.t1592 nfet_06v0 ad=94.5f pd=0.885u as=0.1224p ps=1.04u w=0.36u l=0.6u
X3065 VDD.t2433 a_34124_n12645 a_34036_n12548 VDD.t2432 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3066 VDD.t1641 a_29744_n15604.t17 a_23072_n13432.t6 VDD.t1640 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3067 a_28736_1944 a_22500_n1976 VDD.t1701 VDD.t1700 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3068 a_36700_n18484 a_36612_n18440 VSS.t2966 VSS.t2965 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3069 a_37820_n15348 a_37732_n15304 VSS.t3095 VSS.t3094 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3070 a_39612_n13780 a_39524_n13736 VSS.t2547 VSS.t2546 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3071 a_33686_n11592 a_32854_n12168 a_33538_n12168 VDD.t2859 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3072 a_39612_n10644 a_39524_n10600 VSS.t3923 VSS.t3922 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3073 a_21804_n2273.t1 a_32132_2428 VDD.t3403 VDD.t3402 pfet_06v0 ad=0.5368p pd=3.32u as=0.35315p ps=1.96u w=1.22u l=0.5u
X3074 a_36112_n3456 a_33588_n3461 a_35800_n3456 VSS.t3420 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3075 a_21772_n20836.t0 a_23564_n20836 VSS.t940 VSS.t939 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3076 a_10778_2852.t8 a_10712_4516.t48 VDD.t342 VDD.t341 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3077 VSS.t4304 a_26563_n12212 a_26431_n12168 VSS.t4303 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X3078 a_33086_n12168 a_32650_n12168 a_32854_n12168 VDD.t3186 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X3079 a_27672_n3543 a_27932_n3543 VSS.t3859 VSS.t3858 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X3080 a_13501_n11816.t16 a_13623_n12196.t36 a_11087_n12816.t26 VSS.t1842 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3081 a_44209_1248 a_24481_761.t71 VSS.t809 VSS.t808 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X3082 a_11023_n4162.t4 a_13623_n4162.t30 VSS.t588 VSS.t587 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X3083 a_38268_n9076 a_38180_n9032 VSS.t1667 VSS.t1666 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3084 a_11087_n23528.t18 a_11023_n22908.t32 a_13501_n22528.t14 VDD.t211 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3085 VSS.t1203 a_27190_n5112 a_27666_n5112 VSS.t1202 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X3086 a_35371_n6980 a_28144_n4708 a_22444_n5156 VSS.t3831 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3087 VDD.t4198 a_38380_n9509 a_38292_n9412 VDD.t4197 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3088 VDD.t3436 a_34908_n16916 a_34820_n16872 VDD.t3435 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3089 VDD.t836 a_33776_n5896.t17 a_34708_n5896.t11 VDD.t835 pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3090 a_43756_n5940 a_43668_n5896 VSS.t3652 VSS.t3651 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3091 a_34348_n3140 a_34248_n3310 VDD.t2787 VDD.t2786 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X3092 VSS.t1463 a_26547_n12951 a_26543_n11384 VSS.t1462 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X3093 a_28752_n15348 a_29161_n14476 VDD.t2686 VDD.t2685 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3094 a_32999_n9010 a_32543_n9032 a_32767_n9010 VDD.t3519 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X3095 VDD.t4263 a_47004_n1236 a_46916_n1192 VDD.t2440 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D88 VSS.t4190 a_25940_n17606.t16 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3096 VDD.t1135 a_47452_n12212 a_47364_n12168 VDD.t1134 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3097 a_38256_1564.t5 a_37844_1564 VDD.t4188 VDD.t4187 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3098 VDD.t2656 a_32189_n9860 a_32309_n9240 VDD.t2655 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3099 a_21772_n8292.t1 a_23564_n8292 VSS.t1219 VSS.t1218 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3100 a_21772_n11428.t0 a_23564_n11428 VSS.t1748 VSS.t1747 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3101 VDD.t156 a_26553_377.t5 a_26431_n1192 VDD.t155 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X3102 VDD.t3082 a_45212_n12212 a_45124_n12168 VDD.t3081 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3103 VSS.t164 a_33496_n6659.t27 a_31628_n5940.t4 VSS.t163 nfet_06v0 ad=0.2134p pd=1.85u as=0.1261p ps=1.005u w=0.485u l=0.6u
X3104 a_34908_n20052 a_34820_n20008 VSS.t3954 VSS.t3953 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3105 a_11087_n20850.t23 a_13623_n20230.t34 a_13501_n19850.t13 VSS.t631 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3106 VSS.t3195 a_27055_n1192 a_27531_n617 VSS.t3194 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X3107 VSS.t914 a_21772_n3588.t14 a_13623_n20230.t3 VSS.t913 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3108 a_38403_n799 a_38733_n727 a_38853_n1170 VDD.t1950 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3109 a_11087_n23528.t46 a_2167_3472.t56 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X3110 VDD.t3097 a_29612_n8292 a_28764_n8247 VDD.t3096 pfet_06v0 ad=0.4972p pd=3.14u as=0.4012p ps=1.85u w=1.13u l=0.5u
X3111 VSS.t3172 a_29612_n8292 a_28972_n8247 VSS.t3171 nfet_06v0 ad=0.3586p pd=2.51u as=0.2119p ps=1.335u w=0.815u l=0.6u
X3112 a_13501_n22528.t4 a_13623_n22908.t26 a_11087_n23528.t4 VSS.t221 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3113 a_11087_n23528.t3 a_13623_n22908.t27 a_13501_n22528.t3 VSS.t222 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X3114 a_30532_n8548 a_21916_n6694.t14 a_30348_n8548 VSS.t1100 nfet_06v0 ad=0.1148p pd=1.1u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3115 a_36217_n3500 a_24481_761.t72 VDD.t760 VDD.t759 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X3116 a_25724_n18484 a_25636_n18440 VSS.t2261 VSS.t2260 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3117 a_42116_n1976 a_37859_377 VSS.t2013 VSS.t2012 nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3118 VDD.t678 a_13623_n6840.t34 a_11023_n6840.t13 VDD.t677 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3119 a_44428_n7941 a_44340_n7844 VSS.t1500 VSS.t1499 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3120 VDD.t4229 a_23484_n18917 a_23396_n18820 VDD.t3335 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3121 VSS.t2364 a_30192_n15304.t14 a_24481_761.t4 VSS.t2363 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X3122 a_25831_n11428 a_27526_n9816 VSS.t2471 VSS.t2470 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X3123 VSS.t4310 a_23564_n17700 a_21772_n17700.t2 VSS.t4309 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3124 a_41740_n4805 a_41652_n4708 VSS.t3248 VSS.t3247 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3125 VSS.t2683 a_21692_n13308.t27 a_21604_n13252 VSS.t2682 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3126 a_13623_n9518.t7 a_21772_n17700.t17 VSS.t1049 VSS.t1048 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3127 VSS.t3812 a_23564_n14564.t6 a_21772_n14564.t3 VSS.t3811 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3128 VSS.t2543 a_27820_n16432 a_27192_n14286 VSS.t2542 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X3129 VSS.t4205 a_32108_n2332.t24 a_35156_n325 VSS.t4204 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3130 a_36428_n53 a_36120_n4 VSS.t3062 VSS.t3061 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X3131 VSS.t2685 a_21692_n13308.t28 a_21604_n10116 VSS.t2684 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3132 a_13623_n12196.t4 a_21772_n14564.t13 VSS.t1953 VSS.t1952 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3133 VDD.t3769 a_21692_2431 a_21604_2475 VDD.t3768 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X3134 VSS.t1671 a_21772_n452.t10 a_13623_n22908.t4 VSS.t1670 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3135 VSS.t656 a_29920_n3900.t18 a_33375_n1976 VSS.t655 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X3136 VDD.t1223 a_25612_n6679 a_25524_n6635 VDD.t1222 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X3137 VDD.t3884 a_43980_n6373 a_43892_n6276 VDD.t3883 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3138 VSS.t811 a_24481_761.t73 a_31939_n6976 VSS.t810 nfet_06v0 ad=0.1224p pd=1.04u as=0.134p ps=1.1u w=0.36u l=0.6u
X3139 VDD.t2980 a_42748_n18484 a_42660_n18440 VDD.t2979 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D89 VSS.t525 a_23072_n13432.t72 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3140 a_24716_1208.t1 a_31961_1204 VDD.t3603 VDD.t3602 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3141 VDD.t2818 a_44316_n2804 a_44228_n2760 VDD.t2817 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3142 VDD.t3334 a_43980_n3237 a_43892_n3140 VDD.t3333 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3143 VDD.t98 a_13623_n17552.t34 a_11023_n17552.t14 VDD.t97 pfet_03v3 ad=1.82p pd=6.9u as=0.728p ps=3.32u w=2.8u l=0.28u
X3144 a_30716_n1148 a_30408_n1104 VSS.t3739 VSS.t3738 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X3145 a_23619_n6724 a_23949_n6724 a_24069_n6680 VSS.t987 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X3146 VDD.t33 a_24815_n3588.t15 a_28736_n4633.t1 VDD.t32 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X3147 VDD.t2405 a_40508_n18484 a_40420_n18440 VDD.t2404 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3148 a_11023_n17552.t13 a_13623_n17552.t35 VDD.t100 VDD.t99 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3149 VDD.t762 a_24481_761.t74 a_29744_n15604.t4 VDD.t761 pfet_06v0 ad=0.367p pd=1.92u as=0.2952p ps=1.54u w=0.82u l=0.5u
D90 a_22444_332.t27 VDD.t12 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3150 a_24913_864 a_23136_447 a_24041_816 VSS.t1969 nfet_06v0 ad=93.59999f pd=0.88u as=0.1989p ps=1.465u w=0.36u l=0.6u
X3151 a_23935_n2276 a_23703_n5156.t4 a_23507_n2759 VSS.t3898 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X3152 a_25159_n2276 a_24403_n2414 VSS.t2749 VSS.t2748 nfet_06v0 ad=48.6f pd=0.645u as=0.14985p ps=1.145u w=0.405u l=0.6u
X3153 a_47004_n18484 a_46916_n18440 VSS.t2899 VSS.t2898 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3154 VSS.t1432 a_41392_1944.t18 OUT[4].t5 VSS.t1431 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3155 VDD.t2555 a_35356_n12212 a_35268_n12168 VDD.t2554 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3156 a_47004_n15348 a_46916_n15304 VSS.t4351 VSS.t4350 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3157 a_26103_n1400 a_25647_n1976 VDD.t1926 VDD.t1925 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X3158 VDD.t1238 a_37632_n2020 a_25019_n3588.t1 VDD.t1237 pfet_06v0 ad=0.35315p pd=1.96u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3159 a_29532_n4372.t3 a_29900_n10600.t6 a_29940_n8548 VSS.t3945 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3160 a_44092_n13780 a_44004_n13736 VSS.t3665 VSS.t3664 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3161 VSS.t590 a_13623_n4162.t31 a_2167_3472.t5 VSS.t589 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3162 a_44092_n10644 a_44004_n10600 VSS.t1714 VSS.t1713 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3163 a_11023_n12196.t14 a_13623_n12196.t37 VDD.t1754 VDD.t1753 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3164 a_40060_n18484 a_39972_n18440 VSS.t2901 VSS.t2900 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3165 VSS.t1120 a_25836_n1236.t27 a_30820_n3544 VSS.t1119 nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
D91 VSS.t812 a_24481_761.t75 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3166 a_31788_n5112 a_30452_n5156.t7 a_28736_n4633.t14 VSS.t1081 nfet_06v0 ad=0.1312p pd=1.14u as=0.4161p ps=1.905u w=0.82u l=0.6u
X3167 VDD.t2557 a_23212_n12124 a_23108_n12080 VDD.t2556 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3168 a_40060_n15348 a_39972_n15304 VSS.t4298 VSS.t4297 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3169 VDD.t379 a_10778_2852.t27 a_10712_4516.t23 VDD.t378 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3170 VSS.t407 a_21692_n5468.t26 a_29332_1243 VSS.t406 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3171 a_21772_n3588.t3 a_23564_n3588.t6 VDD.t2917 VDD.t2916 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3172 VDD.t3898 a_29408_1944.t17 OUT[0].t14 VDD.t3897 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3173 a_35916_n12645 a_35828_n12548 VSS.t1864 VSS.t1863 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3174 VDD.t1312 a_13623_n14874.t36 a_11023_n14874.t13 VDD.t1311 pfet_03v3 ad=1.82p pd=6.9u as=0.728p ps=3.32u w=2.8u l=0.28u
X3175 VSS.t3159 a_38984_n1975 a_23564_n452.t0 VSS.t3158 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
D92 VSS.t813 a_24481_761.t76 diode_nd2ps_06v0 pj=1.86u area=0.2052p
D93 VSS.t4191 a_25940_n17606.t17 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3176 a_11023_n14874.t14 a_13623_n14874.t37 VDD.t1314 VDD.t1313 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3177 a_29408_1944.t7 a_22052_1944 VDD.t2718 VDD.t2717 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3178 VDD.t1043 a_30452_n5156.t8 a_28736_n4633.t11 VDD.t1042 pfet_06v0 ad=0.4056p pd=1.805u as=0.2197p ps=1.365u w=0.845u l=0.5u
X3179 a_24233_n5548 a_23072_n13432.t73 VDD.t521 VDD.t520 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X3180 a_24464_n11680 a_22352_n12097 a_24152_n11680 VDD.t1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X3181 a_11087_n18172.t35 a_2167_3472.t75 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X3182 VDD.t1768 a_32579_769 a_28492_332 VDD.t1767 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3183 VSS.t748 a_28156_n6412.t25 a_26440_n5940.t3 VSS.t747 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3184 VDD.t3946 a_40172_n5940 a_40084_n5896 VDD.t3945 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3185 a_13501_n6460.t0 a_13623_n6840.t35 a_11087_n7460.t5 VSS.t738 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3186 VDD.t2325 a_47452_n1236 a_47364_n1192 VDD.t1502 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3187 a_46220_n11077 a_46132_n10980 VSS.t3273 VSS.t3272 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3188 VSS.t563 a_11023_n9518.t31 a_11087_n10138.t11 VSS.t60 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3189 VDD.t3857 a_46332_n20485 a_46244_n20388 VDD.t3856 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3190 a_30901_146 a_30781_n452 VDD.t3323 VDD.t3322 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X3191 a_31461_n7694 a_31341_n8292 VDD.t3974 VDD.t3973 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X3192 VDD.t2471 a_40776_770 a_40672_864 VDD.t2470 pfet_06v0 ad=0.3432p pd=2.44u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3193 a_23527_n2276 a_22164_n2760 VSS.t1947 VSS.t1946 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X3194 a_30095_n13252 a_28940_n2406.t6 a_27820_n16432 VSS.t3082 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X3195 VDD.t3968 a_39612_n7508 a_39524_n7464 VDD.t3967 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3196 a_39724_n15781 a_39636_n15684 VSS.t2119 VSS.t2118 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3197 a_22016_n4257 a_21604_n3844 VSS.t1804 VSS.t1803 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3198 a_31292_n5112 a_24815_n3588.t16 a_28548_n5112 VSS.t24 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3199 a_30092_1564 a_28836_376 VDD.t1612 VDD.t1611 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X3200 VDD.t3208 a_39612_n4372 a_39524_n4328 VDD.t2228 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3201 a_30174_n5112 a_25836_n1236.t28 a_29980_n5112 VSS.t1121 nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X3202 a_31856_n11296 a_29744_n10980 a_31544_n11296 VDD.t3582 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X3203 VDD.t229 a_13623_n22908.t28 a_11023_n22908.t13 VDD.t228 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3204 a_38268_n18484 a_38180_n18440 VSS.t3452 VSS.t3451 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3205 a_26284_1564 a_22096_376 VSS.t4043 VSS.t4042 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3206 a_22568_n1104 a_21604_n708 a_22364_n1104 VSS.t3434 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3207 VDD.t1643 a_29744_n15604.t18 a_23072_n13432.t0 VDD.t1642 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3208 a_26991_860 a_25836_n1236.t29 VSS.t1123 VSS.t1122 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3209 VSS.t1762 a_28009_n12168 a_29360_n12864 VSS.t1761 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3210 a_38268_n15348 a_38180_n15304 VSS.t2541 VSS.t2540 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3211 OUT[3].t4 a_38256_1564.t13 VSS.t180 VSS.t179 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3212 VDD.t907 a_39544_420 a_39352_464 VDD.t906 pfet_06v0 ad=0.2222p pd=1.89u as=0.2424p ps=1.465u w=0.505u l=0.5u
X3213 VSS.t2074 CLK.t10 a_33496_n6659.t6 VSS.t2073 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3214 VDD.t2132 a_39357_n660 a_39477_n1192 VDD.t2131 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3215 a_44876_n17349 a_44788_n17252 VSS.t2335 VSS.t2334 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3216 a_43084_n3237 a_42996_n3140 VSS.t1963 VSS.t1962 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3217 VDD.t3286 a_39556_n4 a_40260_n408 VDD.t3285 pfet_06v0 ad=0.5368p pd=3.32u as=0.3477p ps=1.79u w=1.22u l=0.5u
X3218 VDD.t1087 a_25836_n1236.t30 a_28736_n4633.t8 VDD.t1086 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X3219 a_44876_n7941 a_44788_n7844 VSS.t1020 VSS.t1019 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3220 VDD.t3719 a_39164_n15348 a_39076_n15304 VDD.t3718 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3221 a_44876_n14213 a_44788_n14116 VSS.t2403 VSS.t2402 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3222 VSS.t893 a_4001_4292.t10 a_10778_2852.t13 VSS.t356 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3223 a_26284_1564 a_22096_376 VDD.t3966 VDD.t3965 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X3224 a_44640_1944.t3 a_44004_n1192 VSS.t2578 VSS.t2577 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3225 a_30111_n6221 a_29211_n6724 VSS.t4041 VSS.t4040 nfet_06v0 ad=94.5f pd=0.885u as=0.1224p ps=1.04u w=0.36u l=0.6u
X3226 a_42636_n17349 a_42548_n17252 VSS.t2469 VSS.t2468 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3227 VDD.t820 a_34708_n5896.t25 a_35456_n4628.t5 VDD.t819 pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X3228 a_24200_n14816 a_23360_n15233 a_23912_n15216 VSS.t1513 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3229 a_3935_4156.t0 a_1955_4292.t4 VSS.t1401 VSS.t1400 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X3230 VSS.t4117 a_25685_n7463 a_26095_n7464 VSS.t4116 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X3231 a_11087_n20850.t31 a_2167_3472.t16 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X3232 a_42636_n14213 a_42548_n14116 VSS.t2703 VSS.t2702 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3233 VSS.t592 a_13623_n4162.t32 a_11023_n4162.t3 VSS.t591 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3234 a_13501_n19850.t3 a_11023_n20230.t33 a_11087_n20850.t13 VDD.t1902 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3235 VSS.t2981 a_24041_816 a_23972_864 VSS.t2980 nfet_06v0 ad=93.59999f pd=0.88u as=62.1f ps=0.705u w=0.36u l=0.6u
X3236 VDD.t789 a_28519_n10160.t8 a_28721_n9076.t1 VDD.t788 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3237 a_41392_1944.t1 a_40196_1944 VSS.t3133 VSS.t3132 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3238 a_37484_n11077 a_37396_n10980 VSS.t4011 VSS.t4010 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3239 VSS.t385 a_10778_2852.t28 a_10712_4516.t13 VSS.t384 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3240 a_40260_n408 a_39556_n4 VSS.t3372 VSS.t3371 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3241 a_39357_n5364 a_25020_n8200.t4 VSS.t904 VSS.t903 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3242 VSS.t2995 a_23564_n3588.t7 a_21772_n3588.t2 VSS.t2994 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3243 a_11023_n9518.t3 a_13623_n9518.t26 VSS.t258 VSS.t257 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3244 a_31544_1248 a_29332_1243 a_30604_1515 VDD.t2513 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X3245 VDD.t1993 a_43644_n7508 a_43556_n7464 VDD.t1992 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3246 VDD.t3518 a_32543_n9032 a_32999_n9010 VDD.t3517 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3247 VSS.t260 a_13623_n9518.t27 a_11023_n9518.t2 VSS.t259 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3248 VDD.t3468 a_35356_n20485 a_35268_n20388 VDD.t1461 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3249 a_33533_908 a_24716_1208.t4 VSS.t2271 VSS.t2270 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3250 a_13623_n22908.t5 a_21772_n452.t11 VSS.t1673 VSS.t1672 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3251 VDD.t3874 a_43644_n4372 a_43556_n4328 VDD.t3873 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3252 VDD.t590 a_13623_n20230.t35 a_11023_n20230.t13 VDD.t589 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3253 VDD.t3724 a_33116_n20485 a_33028_n20388 VDD.t2048 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3254 a_28568_n16066 a_28752_n15348 VSS.t3201 VSS.t3200 nfet_06v0 ad=0.1584p pd=1.6u as=0.151p ps=1.185u w=0.36u l=0.6u
X3255 a_24481_761.t5 a_30192_n15304.t15 VSS.t2366 VSS.t2365 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X3256 a_47900_n7508 a_47812_n7464 VSS.t2240 VSS.t2239 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3257 a_33616_n6976 a_24481_761.t77 VSS.t814 VSS.t141 nfet_06v0 ad=43.199997f pd=0.6u as=0.2016p ps=1.48u w=0.36u l=0.6u
X3258 a_27292_n14116 a_27192_n14286 VSS.t2545 VSS.t2544 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3259 VSS.t3596 a_27224_n62 a_27032_51 VSS.t3595 nfet_06v0 ad=0.2016p pd=1.48u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3260 a_31544_n11296 a_29744_n10980 a_30604_n11029 VSS.t3668 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3261 VSS.t65 a_11023_n14874.t32 a_11087_n15494.t24 VSS.t64 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X3262 a_40396_n12645 a_40308_n12548 VSS.t2283 VSS.t2282 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3263 VDD.t2008 a_48012_n15781 a_47924_n15684 VDD.t2007 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3264 a_11087_n15494.t23 a_11023_n14874.t33 VSS.t67 VSS.t66 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3265 a_43420_n2804 a_43332_n2760 VSS.t3857 VSS.t3856 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3266 VDD.t2014 a_46220_n6373 a_46132_n6276 VDD.t2013 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3267 a_31248_n3544 a_25836_n1236.t31 VSS.t1125 VSS.t1124 nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3268 VDD.t660 a_29800_n5940.t17 a_28156_n6412.t10 VDD.t659 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3269 VDD.t3420 a_48012_n12645 a_47924_n12548 VDD.t3419 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3270 VDD.t3465 a_46220_n3237 a_46132_n3140 VDD.t3464 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3271 a_11023_n6840.t14 a_13623_n6840.t36 VDD.t680 VDD.t679 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3272 VSS.t416 a_11023_n17552.t33 a_11087_n18172.t23 VSS.t70 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3273 a_24731_n3124.t0 a_24631_n3588 VDD.t3223 VDD.t3222 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X3274 VDD.t3552 a_33120_n3884 a_33015_n4284 VDD.t3551 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X3275 a_22812_n7376 a_22712_n7420 VSS.t970 VSS.t969 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3276 a_13501_n9138.t13 a_13623_n9518.t28 a_11087_n10138.t20 VSS.t261 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X3277 a_27605_n10600 a_27485_n10068 a_26861_n10135 VDD.t1734 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X3278 a_29856_n1121 a_29444_n708 VSS.t2816 VSS.t2815 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3279 a_30676_n7844 a_30228_n8203 VDD.t3631 VDD.t3630 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X3280 VDD.t1731 a_37820_n12212 a_37732_n12168 VDD.t1730 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3281 a_11087_n18172.t22 a_11023_n17552.t34 VSS.t417 VSS.t72 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X3282 a_22856_n3840 a_22016_n4257 a_22568_n4240 VSS.t3351 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3283 a_27717_n8248 a_27597_n8292 a_26973_n8292 VSS.t2947 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X3284 OUT[0].t13 a_29408_1944.t18 VDD.t3900 VDD.t3899 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3285 VDD.t2030 a_36700_n12212 a_36612_n12168 VDD.t2029 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3286 VDD.t280 a_31548_n10172.t22 a_33588_n3461 VDD.t279 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
D94 a_25940_n17606.t18 VDD.t4120 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3287 VSS.t2345 a_42604_n2020 a_42556_n1976 VSS.t2344 nfet_06v0 ad=0.2132p pd=1.34u as=98.399994f ps=1.06u w=0.82u l=0.6u
X3288 a_25237_n4327 a_24233_n3980 VDD.t1860 VDD.t1859 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3289 a_42748_n12212 a_42660_n12168 VSS.t4070 VSS.t4069 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3290 VSS.t121 a_11023_n12196.t32 a_11087_n12816.t4 VSS.t64 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X3291 a_43084_n15781 a_42996_n15684 VSS.t2064 VSS.t2063 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3292 VSS.t387 a_10778_2852.t29 a_10712_4516.t12 VSS.t386 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3293 a_11087_n12816.t3 a_11023_n12196.t33 VSS.t122 VSS.t66 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3294 a_21892_n12952 a_21772_n12996 VSS.t3725 VSS.t3724 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3295 a_11023_n4162.t15 a_13623_n4162.t33 VDD.t560 VDD.t559 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3296 VDD.t4006 a_46668_n18917 a_46580_n18820 VDD.t4005 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3297 a_32533_n13944 a_32413_n14564 a_31789_n14564 VDD.t1577 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X3298 VDD.t2795 a_39164_n4805 a_39076_n4708 VDD.t2794 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3299 a_40508_n12212 a_40420_n12168 VSS.t3851 VSS.t3850 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3300 VDD.t3869 a_34908_n20052 a_34820_n20008 VDD.t2086 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3301 VDD.t3637 a_41852_n16916 a_41764_n16872 VDD.t3636 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3302 a_34747_952 a_34271_376 VSS.t3531 VSS.t3530 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3303 VDD.t3346 a_41852_n13780 a_41764_n13736 VDD.t3345 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3304 VDD.t2016 a_23816_n3840 a_24233_n3980 VDD.t2015 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X3305 VDD.t2850 a_44428_n18917 a_44340_n18820 VDD.t2849 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3306 a_2167_3472.t6 a_13623_n4162.t34 VSS.t594 VSS.t593 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3307 a_29444_n4328.t3 a_25836_n1236.t32 VDD.t1089 VDD.t1088 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X3308 a_11087_n20850.t40 a_2167_3472.t28 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X3309 a_31787_n3969 a_32359_n4372 VDD.t2525 VDD.t2524 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3310 VDD.t4170 a_39276_n15781 a_39188_n15684 VDD.t4169 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3311 a_10712_4516.t5 a_3935_4156.t10 VSS.t459 VSS.t388 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3312 a_31856_1248 a_29744_1564 a_31544_1248 VDD.t1111 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X3313 a_41616_1564 a_41204_1243 VDD.t1782 VDD.t1781 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X3314 a_41852_n20052 a_41764_n20008 VSS.t2525 VSS.t2524 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3315 a_32104_n3544 a_25836_n1236.t33 VSS.t1127 VSS.t1126 nfet_06v0 ad=0.1722p pd=1.24u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3316 a_21692_n5468.t10 a_26440_n5940.t13 VDD.t355 VDD.t354 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3317 VDD.t4233 a_38156_n12645 a_38068_n12548 VDD.t4232 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3318 VDD.t3645 a_37036_n15781 a_36948_n15684 VDD.t3644 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3319 a_22052_n4708 a_21604_n5067 VSS.t2134 VSS.t2133 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X3320 VSS.t1977 a_11023_n20230.t34 a_11087_n20850.t14 VSS.t54 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3321 a_42448_n1572 a_41684_n1976 a_42244_n1572 VDD.t2384 pfet_06v0 ad=0.4758p pd=2u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3322 a_26981_n8457 a_26861_n8567 VSS.t3003 VSS.t3002 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X3323 a_39612_n18484 a_39524_n18440 VSS.t3039 VSS.t3038 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3324 VDD.t3613 a_31459_n14564 a_30159_n13296 VDD.t3612 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3325 VDD.t3229 a_36520_n3868 a_26388_n17606.t1 VDD.t3228 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3326 a_39612_n15348 a_39524_n15304 VSS.t3741 VSS.t3740 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3327 a_24116_n15216 a_22948_n14820 a_23912_n15216 VDD.t2035 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3328 a_11087_n23528.t22 a_11023_n22908.t33 VSS.t199 VSS.t58 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3329 VDD.t1997 CLK.t11 a_33496_n6659.t3 VDD.t1996 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X3330 VSS.t1785 a_37024_1944.t19 OUT[2].t3 VSS.t1784 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3331 VDD.t452 a_21772_1116.t14 a_13623_n4162.t13 VDD.t451 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3332 a_36744_n1954 a_36388_n1572 VDD.t1030 VDD.t1029 pfet_06v0 ad=0.4488p pd=2.92u as=0.458p ps=2.02u w=1.02u l=0.5u
X3333 a_13501_n14494.t12 a_11023_n14874.t34 a_11087_n15494.t12 VDD.t80 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3334 a_23816_n13248 a_21604_n13252 a_22876_n13692 VDD.t2140 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X3335 VSS.t1434 a_41392_1944.t19 OUT[4].t4 VSS.t1433 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3336 a_28836_376 a_28132_376 VDD.t3695 VDD.t3694 pfet_06v0 ad=0.3477p pd=1.79u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3337 a_21792_n7464 a_21692_n7508.t2 VDD.t4275 VDD.t4274 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3338 a_47116_n7941 a_47028_n7844 VSS.t4333 VSS.t4332 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3339 a_23816_n8544 a_22016_n8961 a_22876_n8988 VSS.t3865 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3340 a_10712_4516.t22 a_10778_2852.t30 VDD.t381 VDD.t380 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3341 VSS.t2600 a_29123_n6679 a_30900_n9032 VSS.t2599 nfet_06v0 ad=0.2911p pd=1.53u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3342 a_23816_n5408 a_22016_n5825 a_22876_n5852 VSS.t3151 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3343 a_39477_n616 a_39357_n660 a_38733_n727 VSS.t2206 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X3344 a_11087_n18172.t12 a_11023_n17552.t35 a_13501_n17172.t12 VDD.t407 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3345 VDD.t1474 a_47004_n5940 a_46916_n5896 VDD.t1473 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3346 VDD.t4204 a_30876_n16916 a_30788_n16872 VDD.t4203 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3347 a_13501_n14494.t7 a_13623_n14874.t38 a_11087_n15494.t7 VSS.t1367 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3348 VSS.t2531 a_26719_n7464 a_27195_n6889 VSS.t2530 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X3349 a_38256_1564.t1 a_37844_1564 VSS.t4262 VSS.t4261 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3350 VDD.t2781 a_47004_n2804 a_46916_n2760 VDD.t2780 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3351 VSS.t1199 a_36217_n3500 a_36112_n3456 VSS.t1198 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X3352 VDD.t662 a_29800_n5940.t18 a_28156_n6412.t9 VDD.t661 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3353 a_34908_n20485 a_34820_n20388 VSS.t1819 VSS.t1818 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3354 VDD.t962 a_37820_n20485 a_37732_n20388 VDD.t961 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3355 a_10712_4516.t6 a_3935_4156.t11 VSS.t460 VSS.t390 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3356 VSS.t995 a_23887_n5156 a_23823_n5111 VSS.t994 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X3357 a_38403_n799 a_38733_n727 a_38853_n617 VSS.t2025 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X3358 VDD.t3075 a_47004_n12212 a_46916_n12168 VDD.t3074 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3359 VDD.t2635 a_26328_n6654.t19 a_21692_n13308.t10 VDD.t2634 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3360 a_31685_n9816 a_31565_n9860 VSS.t2292 VSS.t2291 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X3361 a_13501_n11816.t2 a_11023_n12196.t34 a_11087_n12816.t12 VDD.t134 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3362 a_25769_860 a_24481_761.t78 a_25137_864 VSS.t815 nfet_06v0 ad=48.6f pd=0.645u as=0.3123p ps=2.38u w=0.405u l=0.6u
D95 VSS.t816 a_24481_761.t79 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3363 a_47004_n9076 a_46916_n9032 VSS.t2101 VSS.t2100 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3364 a_30876_n20052 a_30788_n20008 VSS.t2140 VSS.t2139 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3365 a_31664_n13292 a_31548_n10172.t23 VDD.t282 VDD.t281 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X3366 a_28004_860 a_27884_332.t4 VSS.t754 VSS.t753 nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3367 a_25685_n7463 a_24681_n7116 VDD.t3193 VDD.t3192 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3368 VDD.t4239 a_40060_n12212 a_39972_n12168 VDD.t4238 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3369 a_29408_1944.t6 a_22052_1944 VDD.t2716 VDD.t2715 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
D96 CLK.t12 VDD.t1998 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3370 a_43980_n12645 a_43892_n12548 VSS.t3044 VSS.t3043 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D97 a_21804_n2273.t11 VDD.t1268 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3371 VSS.t4035 a_31235_n9860 a_29992_n11150 VSS.t4034 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3372 VSS.t1472 a_31760_n12168 a_33280_n13248 VSS.t1471 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3373 a_23136_447 a_22724_860.t4 VSS.t917 VSS.t916 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3374 VDD.t2664 a_45660_332 a_45572_376 VDD.t2663 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3375 a_13501_n11816.t17 a_13623_n12196.t38 a_11087_n12816.t27 VSS.t1843 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3376 a_13623_n14874.t13 a_21772_n11428.t18 VDD.t306 VDD.t305 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3377 a_41740_n12645 a_41652_n12548 VSS.t3244 VSS.t3243 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3378 a_11087_n18172.t3 a_13623_n17552.t36 a_13501_n17172.t3 VSS.t94 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3379 a_41740_n9509 a_41652_n9412 VSS.t2719 VSS.t2718 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3380 a_21692_n18484 a_21604_n18440 VSS.t3058 VSS.t3057 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3381 VSS.t12 a_22444_332.t28 a_29659_n14820 VSS.t11 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3382 a_29956_n2760 a_24815_n3588.t17 a_29732_n2760 VDD.t34 pfet_06v0 ad=0.3172p pd=1.74u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3383 a_24481_761.t6 a_30192_n15304.t16 VSS.t2368 VSS.t2367 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X3384 VDD.t1545 a_34403_332 a_34271_376 VDD.t1544 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X3385 a_21692_n15348 a_21604_n15304 VSS.t2056 VSS.t2055 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3386 VDD.t2137 a_23324_n7420 a_23220_n7376 VDD.t2136 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3387 VDD.t3344 a_23036_n18917 a_22948_n18820 VDD.t3343 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3388 VSS.t2370 a_30192_n15304.t17 a_24481_761.t7 VSS.t2369 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X3389 VSS.t424 a_28721_n9076.t8 a_30136_n10600 VSS.t423 nfet_06v0 ad=0.218p pd=1.52u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3390 VDD.t4277 a_46668_n9509 a_46580_n9412 VDD.t4276 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3391 a_26755_n16132 a_27085_n16132 a_27205_n16088 VSS.t1958 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X3392 VDD.t4223 a_24578_n2020 a_24698_n1400 VDD.t4222 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3393 a_23228_n6679 a_23479_n5156 a_23415_n5111 VSS.t2314 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X3394 a_26776_1248 a_25936_1564 a_26488_1564 VSS.t1486 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3395 VDD.t1416 a_39164_n9076 a_39076_n9032 VDD.t1415 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3396 a_13501_n22528.t13 a_11023_n22908.t34 a_11087_n23528.t17 VDD.t212 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3397 VDD.t1359 a_38604_n7941 a_38516_n7844 VDD.t1358 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3398 VDD.t194 a_38256_1564.t14 OUT[3].t13 VDD.t193 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3399 a_21692_n5468.t9 a_26440_n5940.t14 VDD.t320 VDD.t319 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3400 VSS.t1258 a_38403_n5503 a_36773_n5468 VSS.t1257 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3401 a_30808_n10116 a_30136_n10600 VSS.t1264 VSS.t1263 nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X3402 a_11087_n23528.t16 a_11023_n22908.t35 a_13501_n22528.t12 VDD.t213 pfet_03v3 ad=0.728p pd=3.32u as=1.82p ps=6.9u w=2.8u l=0.28u
D98 VSS.t526 a_23072_n13432.t74 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3403 a_37024_1944.t0 a_36388_1944 VSS.t1736 VSS.t1735 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3404 VDD.t1045 a_30452_n5156.t9 a_27259_804.t1 VDD.t1044 pfet_06v0 ad=0.5368p pd=3.32u as=0.4575p ps=1.97u w=1.22u l=0.5u
X3405 a_37605_n3544 a_22052_n4708 VSS.t3697 VSS.t3696 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3406 VDD.t3291 a_38268_n12212 a_38180_n12168 VDD.t3290 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3407 a_44092_n18484 a_44004_n18440 VSS.t3033 VSS.t3032 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3408 VDD.t2018 a_26844_n20485 a_26756_n20388 VDD.t2017 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3409 a_29295_n1400 a_28671_n1976 a_29127_n1400 VDD.t3782 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3410 VDD.t1098 a_43980_n17349 a_43892_n17252 VDD.t1097 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3411 a_44092_n15348 a_44004_n15304 VSS.t2147 VSS.t2146 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3412 a_43416_1248 a_41616_1564 a_42476_1515 VSS.t2821 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3413 a_39948_n12645 a_39860_n12548 VSS.t980 VSS.t979 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3414 VDD.t1246 a_43980_n14213 a_43892_n14116 VDD.t1245 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3415 a_31451_n7508 a_31799_n7508 VDD.t1551 VDD.t1550 pfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X3416 VDD.t1764 a_24604_n20485 a_24516_n20388 VDD.t1763 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3417 VDD.t1248 a_41740_n17349 a_41652_n17252 VDD.t1247 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3418 VSS.t1154 a_21916_n1975 a_21828_n1931 VSS.t1153 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3419 a_37708_n12645 a_37620_n12548 VSS.t1028 VSS.t1027 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3420 a_28156_n6412.t8 a_29800_n5940.t19 VDD.t664 VDD.t663 pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3421 a_47564_n7941 a_47476_n7844 VSS.t2382 VSS.t2381 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3422 a_30787_n12167 a_27988_n4328 a_30599_n12167 VDD.t1512 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3423 VDD.t1250 a_40620_n17349 a_40532_n17252 VDD.t1249 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3424 VDD.t1252 a_41740_n14213 a_41652_n14116 VDD.t1251 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3425 a_33672_n10112 a_31872_n10529 a_32732_n10556 VSS.t3822 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3426 VSS.t934 a_32413_n12996 a_32533_n12952 VSS.t933 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3427 VDD.t1371 a_40620_n14213 a_40532_n14116 VDD.t1370 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3428 VDD.t1273 a_33252_n1192 a_29900_760.t1 VDD.t1272 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3429 a_21916_n1975 a_25836_n1236.t34 VSS.t1129 VSS.t1128 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X3430 VDD.t1165 a_25237_n4327 a_25759_n3544 VDD.t1164 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X3431 VDD.t4091 a_35456_n4628.t19 a_32108_n2332.t10 VDD.t4090 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3432 a_36364_n7941 a_36276_n7844 VSS.t2485 VSS.t2484 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3433 a_11087_n23528.t47 a_2167_3472.t55 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X3434 a_30584_n1954 a_29444_n4328.t8 VSS.t1563 VSS.t1562 nfet_06v0 ad=0.1584p pd=1.6u as=0.151p ps=1.185u w=0.36u l=0.6u
X3435 VDD.t1890 a_39500_n12645 a_39412_n12548 VDD.t1889 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3436 VDD.t4212 a_47452_n5940 a_47364_n5896 VDD.t4211 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3437 a_31628_n5940.t23 a_33496_n6659.t28 VDD.t174 VDD.t173 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3438 a_39500_n6373 a_39412_n6276 VSS.t2358 VSS.t2357 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3439 VSS.t528 a_23072_n13432.t75 a_23024_n13248 VSS.t527 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3440 VDD.t3579 a_47452_n2804 a_47364_n2760 VDD.t3578 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3441 a_48012_n11077 a_47924_n10980 VSS.t3060 VSS.t3059 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3442 a_27932_n3543 a_23703_n5156.t5 a_28433_n3844 VSS.t3899 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X3443 a_37372_n7508 a_37284_n7464 VSS.t4076 VSS.t4075 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3444 a_13501_n9138.t5 a_11023_n9518.t32 a_11087_n10138.t12 VDD.t546 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3445 VDD.t974 a_34232_n2272 a_34649_n2412 VDD.t973 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3446 VSS.t2763 a_11023_n4162.t33 a_2167_3472.t36 VDD.t2696 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3447 a_24752_n8292 a_25020_n8200.t5 VDD.t845 VDD.t844 pfet_06v0 ad=0.2486p pd=2.01u as=0.35315p ps=1.96u w=0.565u l=0.5u
X3448 VDD.t3109 a_43196_n9076 a_43108_n9032 VDD.t3108 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3449 VSS.t1801 a_42157_n660 a_42277_n616 VSS.t1800 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3450 VDD.t4106 a_42636_n7941 a_42548_n7844 VDD.t4105 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3451 VDD.t3566 a_41180_n20485 a_41092_n20388 VDD.t3565 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3452 OUT[3].t3 a_38256_1564.t15 VSS.t182 VSS.t181 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3453 a_35692_n15781 a_35604_n15684 VSS.t2463 VSS.t2462 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3454 a_30684_860 a_29900_760.t15 a_30372_376 VSS.t2302 nfet_06v0 ad=98.399994f pd=1.06u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3455 a_30662_n3844 a_29920_n3900.t19 a_30468_n3844 VSS.t657 nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X3456 VDD.t2540 a_42636_n4805 a_42548_n4708 VDD.t2539 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3457 VDD.t3564 a_40060_n20485 a_39972_n20388 VDD.t3563 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3458 OUT[0].t12 a_29408_1944.t19 VDD.t3902 VDD.t3901 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3459 a_47452_n9076 a_47364_n9032 VSS.t2198 VSS.t2197 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3460 a_11023_n12196.t15 a_13623_n12196.t39 VDD.t1756 VDD.t1755 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3461 a_33452_n15781 a_33364_n15684 VSS.t4078 VSS.t4077 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3462 a_25899_n3752 a_25423_n4328 VSS.t1391 VSS.t1390 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3463 VDD.t1145 a_39357_n5364 a_39477_n5896 VDD.t1144 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3464 a_25685_n7463 a_24681_n7116 VSS.t3280 VSS.t3279 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X3465 VDD.t86 a_21772_n8292.t19 a_13623_n17552.t10 VDD.t85 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3466 VDD.t3374 a_38828_n17349 a_38740_n17252 VDD.t3373 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3467 a_13501_n6460.t8 a_11023_n6840.t33 a_11087_n7460.t22 VDD.t114 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3468 a_28232_n12606 a_27639_n12537 a_28968_n12864 VSS.t2155 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3469 VDD.t2762 a_39357_n2228 a_39477_n2760 VDD.t2761 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3470 a_46668_n17349 a_46580_n17252 VSS.t4232 VSS.t4231 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3471 VSS.t2495 a_22668_n14864.t3 a_22264_n8988 VSS.t1952 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X3472 VDD.t3378 a_38828_n14213 a_38740_n14116 VDD.t3377 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3473 VDD.t3577 a_45212_n9076 a_45124_n9032 VDD.t3576 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3474 a_33776_n5896.t2 a_31628_n5940.t40 VSS.t136 VSS.t135 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3475 a_46668_n14213 a_46580_n14116 VSS.t2449 VSS.t2448 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3476 a_34708_n5896.t10 a_33776_n5896.t18 VDD.t838 VDD.t837 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3477 a_44428_n17349 a_44340_n17252 VSS.t4252 VSS.t4251 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3478 a_40396_n7941 a_40308_n7844 VSS.t2727 VSS.t2726 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3479 a_22364_n8944 a_22264_n8988 VSS.t2997 VSS.t2996 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3480 VDD.t3380 a_30764_n17349 a_30676_n17252 VDD.t3379 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3481 a_23816_n10112 a_22016_n10529 a_22876_n10556 VSS.t1954 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3482 a_44428_n14213 a_44340_n14116 VSS.t4240 VSS.t4239 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3483 VSS.t461 a_3935_4156.t12 a_10712_4516.t7 VSS.t372 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3484 a_22364_n5808 a_22264_n5852 VSS.t1585 VSS.t1584 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3485 a_31628_n5940.t3 a_33496_n6659.t29 VSS.t166 VSS.t165 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X3486 VDD.t2765 a_43644_n705 a_43556_n661 VDD.t2764 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X3487 a_43532_n6373 a_43444_n6276 VSS.t4228 VSS.t4227 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3488 VDD.t3296 a_43868_n1669 a_43780_n1572 VDD.t3295 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3489 a_39276_n11077 a_39188_n10980 VSS.t2937 VSS.t2936 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3490 VDD.t2600 a_25544_n16412 a_23564_n11428 VDD.t2599 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3491 VDD.t1440 a_40956_n10644 a_40868_n10600 VDD.t1439 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3492 a_27531_n617 a_27055_n1192 a_27279_n1170 VSS.t3193 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
D99 a_23072_n13432.t76 VDD.t522 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3493 VDD.t2012 a_n263_3472.t18 a_137_4292 VDD.t2011 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X3494 a_28225_n4327 a_22164_n2760 a_27932_n3543 VDD.t1870 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3495 a_11023_n6840.t15 a_13623_n6840.t37 VDD.t682 VDD.t681 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3496 a_37036_n11077 a_36948_n10980 VSS.t3288 VSS.t3287 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3497 VDD.t3012 a_38268_n20485 a_38180_n20388 VDD.t3011 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3498 VDD.t4161 a_41852_n20052 a_41764_n20008 VDD.t4160 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3499 a_26553_377.t0 a_25817_804 VSS.t3220 VSS.t3219 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X3500 VDD.t2605 a_21692_n5111.t4 a_21604_n5067 VDD.t398 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X3501 a_11087_n10138.t13 a_11023_n9518.t33 VSS.t564 VSS.t62 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3502 a_28736_n4633.t5 a_21916_n6694.t15 VDD.t1061 VDD.t1060 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X3503 VDD.t3759 a_25237_n5895 a_25530_n5112 VDD.t3758 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X3504 a_23472_n6976 a_23324_n7420 a_23304_n6976 VSS.t2215 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3505 a_40956_n16916 a_40868_n16872 VSS.t4337 VSS.t4336 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3506 VDD.t3385 a_37932_n9509 a_37844_n9412 VDD.t3384 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3507 VSS.t3701 a_34649_n2412 a_34544_n2272 VSS.t3700 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X3508 a_21692_n5468.t3 a_26440_n5940.t15 VSS.t332 VSS.t331 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X3509 VDD.t840 a_33776_n5896.t19 a_34708_n5896.t9 VDD.t839 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3510 VSS.t110 a_11023_n6840.t34 a_11087_n7460.t13 VSS.t70 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3511 VSS.t1710 a_30555_n13780 a_28927_n10160 VSS.t1709 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X3512 VSS.t1787 a_37024_1944.t20 OUT[2].t2 VSS.t1786 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3513 a_30740_n7464 a_30036_n7464 VDD.t3065 VDD.t3064 pfet_06v0 ad=0.3477p pd=1.79u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3514 VDD.t266 a_13623_n9518.t29 a_11023_n9518.t13 VDD.t265 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3515 a_42188_n12645 a_42100_n12548 VSS.t3645 VSS.t3644 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3516 a_38380_n18917 a_38292_n18820 VSS.t3250 VSS.t3249 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3517 a_35456_n4628.t0 a_34708_n5896.t26 VSS.t870 VSS.t869 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3518 a_11087_n23528.t48 a_2167_3472.t54 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
D100 a_21692_n6694.t21 VDD.t641 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3519 VSS.t2187 a_43725_908 a_43845_952 VSS.t2186 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3520 a_11023_n4162.t14 a_13623_n4162.t35 VDD.t562 VDD.t561 pfet_03v3 ad=0.728p pd=3.32u as=1.82p ps=6.9u w=2.8u l=0.28u
X3521 VDD.t4093 a_35456_n4628.t20 a_32108_n2332.t9 VDD.t4092 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3522 a_46108_n5940 a_46020_n5896 VSS.t1659 VSS.t1658 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3523 a_11087_n15494.t32 a_2167_3472.t11 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X3524 a_36140_n18917 a_36052_n18820 VSS.t3246 VSS.t3245 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3525 a_31628_n5940.t22 a_33496_n6659.t30 VDD.t176 VDD.t175 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3526 a_38380_n9509 a_38292_n9412 VSS.t4272 VSS.t4271 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3527 VSS.t740 a_13623_n6840.t38 a_11023_n6840.t16 VSS.t739 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X3528 a_22444_n5156 a_28144_n4708 VDD.t3756 VDD.t3755 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X3529 a_2167_3472.t7 a_13623_n4162.t36 VSS.t596 VSS.t595 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3530 a_31032_n10116 a_28721_n9076.t9 a_30808_n10116 VSS.t425 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3531 a_34162_n11593 a_33686_n11592 a_33910_n12146 VSS.t3155 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X3532 a_27225_n1572.t1 a_26495_n1976 VDD.t2390 VDD.t2389 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X3533 a_25600_n5895 a_24672_n11339 a_25412_n5895 VDD.t1891 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3534 a_42300_n9076 a_42212_n9032 VSS.t2457 VSS.t2456 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3535 VDD.t2824 a_39612_n12212 a_39524_n12168 VDD.t2823 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3536 a_28225_n4327 a_23703_n5156.t6 VDD.t3818 VDD.t3817 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3537 a_33776_n5896.t4 a_31628_n5940.t41 VDD.t150 VDD.t149 pfet_06v0 ad=0.2952p pd=1.54u as=0.3608p ps=2.52u w=0.82u l=0.5u
X3538 VSS.t1436 a_41392_1944.t20 OUT[4].t3 VSS.t1435 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3539 a_28736_n4633.t9 a_25836_n1236.t35 VDD.t1091 VDD.t1090 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X3540 a_11087_n20850.t15 a_11023_n20230.t35 a_13501_n19850.t2 VDD.t1903 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3541 VDD.t1957 a_23542_n1754 a_23642_n1400 VDD.t1956 pfet_06v0 ad=0.1656p pd=1.28u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3542 VDD.t1476 a_34392_n9815 a_28335_n10644 VDD.t1475 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
D101 VSS.t234 a_26388_n17606.t9 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3543 a_28529_1248 a_24481_761.t80 VSS.t818 VSS.t817 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X3544 a_42372_1564 a_24481_761.t81 VDD.t764 VDD.t763 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X3545 VSS.t3956 a_38403_n799 a_33820_n452.t0 VSS.t3955 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3546 VDD.t1290 a_43644_n16916 a_43556_n16872 VDD.t1289 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3547 a_11087_n7460.t6 a_13623_n6840.t39 a_13501_n6460.t5 VSS.t741 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X3548 VSS.t3743 a_23564_n452.t4 a_21772_n452.t2 VSS.t3742 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3549 VDD.t2724 a_25076_n4.t3 a_32132_n4708 VDD.t2723 pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X3550 VDD.t2070 a_30876_n20052 a_30788_n20008 VDD.t2069 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3551 VDD.t3689 a_43644_n13780 a_43556_n13736 VDD.t3688 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3552 a_25132_n16432 a_25831_n12996 a_25767_n12951 VSS.t2612 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X3553 a_42972_n20485 a_42884_n20388 VSS.t2341 VSS.t2340 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3554 a_32482_n12168 a_32026_n12168 VDD.t3704 VDD.t3703 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X3555 VDD.t1180 a_41404_n16916 a_41316_n16872 VDD.t1179 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3556 a_28153_1204 a_27736_1248 a_28529_1248 VSS.t3461 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X3557 VDD.t1292 a_45660_n9076 a_45572_n9032 VDD.t1291 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3558 a_22904_n12080 a_21940_n11684 a_22700_n12080 VSS.t2274 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3559 a_31459_n12996 a_31789_n12996 a_31909_n12398 VDD.t4299 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3560 VDD.t934 a_42188_n17349 a_42100_n17252 VDD.t933 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3561 VDD.t3092 a_41404_n13780 a_41316_n13736 VDD.t3091 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3562 VSS.t633 a_13623_n20230.t36 a_11023_n20230.t3 VSS.t632 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3563 VDD.t1298 a_42188_n14213 a_42100_n14116 VDD.t1297 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3564 a_30452_n5156.t2 a_36744_n1954 VDD.t2806 VDD.t2805 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3565 a_40732_n20485 a_40644_n20388 VSS.t2465 VSS.t2464 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3566 a_13623_n17552.t9 a_21772_n8292.t20 VDD.t68 VDD.t67 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3567 a_11023_n20230.t2 a_13623_n20230.t37 VSS.t635 VSS.t634 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X3568 a_33120_n3884 a_32108_n2332.t25 VSS.t4207 VSS.t4206 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3569 a_43644_n20052 a_43556_n20008 VSS.t1239 VSS.t1238 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3570 VDD.t3167 a_34908_n18484 a_34820_n18440 VDD.t3166 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3571 a_25076_n4.t0 a_24628_n363 VSS.t1981 VSS.t1980 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X3572 a_32432_n2689 a_32020_n2276 VSS.t3108 VSS.t3107 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3573 VSS.t4193 a_25940_n17606.t19 a_35371_n6980 VSS.t4192 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3574 a_31043_n13248 a_30903_n13780 a_30555_n13780 VSS.t2579 nfet_06v0 ad=0.134p pd=1.1u as=0.176p ps=1.68u w=0.4u l=0.6u
X3575 a_43980_n6373 a_43892_n6276 VSS.t3968 VSS.t3967 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3576 VSS.t224 a_13623_n22908.t29 a_11023_n22908.t2 VSS.t223 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3577 a_13623_n6840.t11 a_21772_n20836.t20 VDD.t628 VDD.t627 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3578 VSS.t69 a_11023_n14874.t35 a_11087_n15494.t22 VSS.t68 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3579 a_46668_n4805 a_46580_n4708 VSS.t2210 VSS.t2209 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3580 a_22856_n13248 a_22016_n13665 a_22568_n13648 VSS.t3926 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3581 a_41404_n20052 a_41316_n20008 VSS.t1343 VSS.t1342 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3582 VDD.t614 a_29920_n3900.t20 a_22444_332.t2 VDD.t613 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3583 a_28736_n4633.t6 a_21916_n6694.t16 VDD.t1063 VDD.t1062 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X3584 VDD.t524 a_23072_n13432.t77 a_29211_n6724 VDD.t523 pfet_06v0 ad=0.29465p pd=1.74u as=0.26p ps=1.52u w=1u l=0.5u
X3585 a_25137_864 a_24481_761.t82 VDD.t766 VDD.t765 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X3586 VSS.t2473 a_24760_n11383 a_24672_n11339 VSS.t2472 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X3587 VSS.t1102 a_21916_n6694.t17 a_24180_n5112 VSS.t1101 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3588 a_11087_n10138.t14 a_11023_n9518.t34 a_13501_n9138.t6 VDD.t547 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3589 a_22116_n9412 a_21996_n12996.t11 a_21872_n9394 VDD.t3489 pfet_06v0 ad=0.3172p pd=1.74u as=0.4248p ps=1.94u w=1.22u l=0.5u
X3590 VDD.t3289 a_27302_n9816 a_27758_n9262 VDD.t1930 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3591 a_11087_n23528.t49 a_2167_3472.t53 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X3592 a_34460_n18484 a_34372_n18440 VSS.t3286 VSS.t3285 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3593 a_34428_n452.t1 a_37785_n364 VDD.t1827 VDD.t1826 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3594 VSS.t168 a_33496_n6659.t31 a_31628_n5940.t2 VSS.t167 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X3595 VSS.t689 a_21692_n6694.t22 a_29540_n11728 VSS.t688 nfet_06v0 ad=0.104p pd=0.92u as=0.14p ps=1.1u w=0.4u l=0.6u
X3596 a_37372_n13780 a_37284_n13736 VSS.t4121 VSS.t4120 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3597 a_2167_3472.t37 a_11023_n4162.t34 VSS.t2764 VDD.t2697 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3598 a_37372_n10644 a_37284_n10600 VSS.t1894 VSS.t1893 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3599 VSS.t418 a_11023_n17552.t36 a_11087_n18172.t21 VSS.t54 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3600 a_35800_n3456 a_34000_n3140 a_34860_n3189 VSS.t2775 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3601 VSS.t51 a_21772_n8292.t21 a_13623_n17552.t1 VSS.t50 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3602 a_32395_n8456 a_31919_n9032 VSS.t2222 VSS.t2221 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3603 a_13501_n9138.t12 a_13623_n9518.t30 a_11087_n10138.t29 VSS.t262 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3604 a_32220_n18484 a_32132_n18440 VSS.t2285 VSS.t2284 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3605 a_31548_n10172.t1 a_33496_n8222.t19 VSS.t304 VSS.t303 nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X3606 VSS.t3331 a_27628_n3841 a_27540_n3797 VSS.t3330 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
D102 VSS.t529 a_23072_n13432.t78 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3607 VDD.t2961 a_42860_n101 a_42772_n4 VDD.t2960 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3608 VSS.t123 a_11023_n12196.t35 a_11087_n12816.t2 VSS.t68 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3609 VDD.t915 a_32668_n16916 a_32580_n16872 VDD.t914 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3610 a_24964_n14116 a_24516_n14475 VSS.t4058 VSS.t4057 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X3611 a_25084_1564 a_24628_1252 VSS.t3717 VSS.t3716 nfet_06v0 ad=0.3608p pd=2.52u as=0.2344p ps=1.56u w=0.82u l=0.6u
X3612 VSS.t4296 a_26499_n2732 a_26495_n2272 VSS.t4295 nfet_06v0 ad=93.59999f pd=0.88u as=86.399994f ps=0.84u w=0.36u l=0.6u
X3613 VSS.t1532 a_34392_n9815 a_28335_n10644 VSS.t1531 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X3614 a_11087_n20850.t38 a_2167_3472.t25 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X3615 VSS.t2242 a_42771_769 a_40776_770 VSS.t2241 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3616 a_46556_n5940 a_46468_n5896 VSS.t4331 VSS.t4330 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3617 a_11087_n23528.t50 a_2167_3472.t52 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X3618 a_31996_n20485 a_31908_n20388 VSS.t2475 VSS.t2474 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3619 VDD.t960 a_30428_n16916 a_30340_n16872 VDD.t959 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D103 VSS.t819 a_24481_761.t83 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3620 VDD.t2195 a_46108_n1669 a_46020_n1572 VDD.t2194 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3621 a_13623_n20230.t2 a_21772_n3588.t15 VSS.t906 VSS.t905 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3622 a_33672_n10112 a_31460_n10116 a_32732_n10556 VDD.t1278 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X3623 VSS.t462 a_3935_4156.t13 a_10712_4516.t8 VSS.t374 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X3624 VDD.t3168 a_39612_n20485 a_39524_n20388 VDD.t2044 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3625 a_38403_n2367 a_38733_n2295 a_38853_n2185 VSS.t2823 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X3626 VDD.t1202 a_34796_n15348 a_34708_n15304 VDD.t1201 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3627 VDD.t3197 a_44540_332 a_44452_376 VDD.t3196 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3628 a_32073_n844 a_31656_n704 a_32449_n704 VSS.t2450 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X3629 VDD.t3319 a_44092_n12212 a_44004_n12168 VDD.t3318 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3630 a_32668_n20052 a_32580_n20008 VSS.t1461 VSS.t1460 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3631 a_36388_1944 a_35940_2475 VDD.t3438 VDD.t3437 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X3632 a_40859_2428 a_27884_332.t5 a_21996_332.t0 VSS.t710 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3633 a_23981_464 a_22724_860.t5 a_23728_464 VDD.t861 pfet_06v0 ad=0.101p pd=0.905u as=0.19315p ps=1.27u w=0.505u l=0.5u
X3634 a_13623_n22908.t4 a_21772_n452.t12 VSS.t1675 VSS.t1674 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3635 VDD.t178 a_33496_n6659.t32 a_31628_n5940.t21 VDD.t177 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3636 VSS.t531 a_23072_n13432.t79 a_24368_n14816 VSS.t530 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3637 a_45772_n12645 a_45684_n12548 VSS.t961 VSS.t960 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3638 VDD.t2893 a_22876_n1148 a_22772_n1104 VDD.t2892 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3639 a_23619_n12996 a_23949_n12996 a_24069_n12952 VSS.t1248 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X3640 a_30428_n20052 a_30340_n20008 VSS.t1465 VSS.t1464 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3641 a_13501_n14494.t11 a_11023_n14874.t36 a_11087_n15494.t11 VDD.t81 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3642 a_31412_n2276 a_24631_n3588 a_31392_n2760 VSS.t3310 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3643 a_42636_n3237 a_42548_n3140 VSS.t3606 VSS.t3605 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3644 a_23024_n10112 a_22876_n10556 a_22856_n10112 VSS.t1168 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3645 a_21772_n11428.t5 a_23564_n11428 VDD.t1667 VDD.t1666 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3646 a_43532_n12645 a_43444_n12548 VSS.t2511 VSS.t2510 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3647 a_26590_n4536 a_26154_n4536 a_26358_n4618 VDD.t1884 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X3648 VSS.t2687 a_21692_n13308.t29 a_21940_n11684 VSS.t2686 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3649 VDD.t3084 a_30451_n452 a_28456_n364 VDD.t3083 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3650 VDD.t308 a_21772_n11428.t19 a_13623_n14874.t12 VDD.t307 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3651 a_23484_n18484 a_23396_n18440 VSS.t2388 VSS.t2387 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3652 OUT[4].t2 a_41392_1944.t21 VSS.t1438 VSS.t1437 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3653 a_39052_n7941 a_38964_n7844 VSS.t4150 VSS.t4149 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3654 a_34652_n11391 a_34089_n10252 VSS.t1579 VSS.t1578 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X3655 VDD.t2775 a_44876_n11077 a_44788_n10980 VDD.t2774 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3656 VSS.t3376 a_27302_n9816 a_27778_n9816 VSS.t3375 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
D104 VSS.t532 a_23072_n13432.t80 diode_nd2ps_06v0 pj=1.86u area=0.2052p
D105 VSS.t4139 a_22140_n6694.t14 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3657 VDD.t2565 a_28744_n14432 a_29161_n14476 VDD.t2564 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X3658 a_31628_n5940.t20 a_33496_n6659.t33 VDD.t180 VDD.t179 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3659 a_23324_n7420 a_23016_n7376 VSS.t1558 VSS.t1557 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X3660 a_45648_1564.t2 a_40652_n1572 VSS.t925 VSS.t924 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3661 VDD.t14 a_22444_332.t29 a_21996_332.t1 VDD.t13 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X3662 a_31961_1204 a_24481_761.t84 VDD.t768 VDD.t767 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X3663 a_22364_n1104 a_22264_n1148.t3 VSS.t3785 VSS.t3784 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3664 VDD.t4043 a_42636_n11077 a_42548_n10980 VDD.t4042 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3665 a_21772_n8292.t4 a_23564_n8292 VDD.t1172 VDD.t1171 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3666 OUT[0].t11 a_29408_1944.t20 VDD.t3904 VDD.t3903 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3667 VSS.t184 a_38256_1564.t16 OUT[3].t2 VSS.t183 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3668 VDD.t3728 a_25836_n1236.t36 a_22444_332.t1 VDD.t3727 pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3669 a_24074_n1976 a_23954_n2020 VSS.t2281 VSS.t2280 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3670 VDD.t564 a_13623_n4162.t37 a_11023_n4162.t13 VDD.t563 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3671 VDD.t1410 a_42188_n9509 a_42100_n9412 VDD.t1409 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3672 a_31960_n13648 a_31559_n13692 a_30903_n13780 VSS.t4073 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3673 a_13501_n11816.t1 a_11023_n12196.t36 a_11087_n12816.t11 VDD.t135 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3674 VDD.t1219 a_22140_n15348 a_22052_n15304 VDD.t1218 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3675 VDD.t1412 a_45324_n7941 a_45236_n7844 VDD.t1411 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3676 a_11087_n18172.t11 a_11023_n17552.t37 a_13501_n17172.t11 VDD.t408 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3677 a_46220_n15781 a_46132_n15684 VSS.t1144 VSS.t1143 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3678 VDD.t2773 a_29756_n20485 a_29668_n20388 VDD.t2772 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3679 VDD.t1017 a_21772_n17700.t18 a_13623_n9518.t6 VDD.t1016 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3680 a_27259_804.t1 a_30452_n5156.t10 VDD.t1047 VDD.t1046 pfet_06v0 ad=0.4575p pd=1.97u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3681 a_31292_n2804 a_31324_n4372 VSS.t4101 VSS.t4100 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X3682 VDD.t3203 a_45324_n4805 a_45236_n4708 VDD.t3202 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3683 VSS.t3588 a_35064_n11383 a_28300_n15348 VSS.t3587 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X3684 a_21692_2431 a_28153_1204 VDD.t3432 VDD.t3431 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3685 a_22568_n1104 a_22016_n1121 a_22364_n1104 VDD.t3361 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3686 a_13623_n9518.t4 a_21772_n17700.t19 VDD.t1019 VDD.t1018 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3687 VDD.t1876 a_21772_n14564.t14 a_13623_n12196.t9 VDD.t1875 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3688 VSS.t3867 a_29800_n9815 a_22220_n12996 VSS.t2038 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X3689 VDD.t2415 a_43980_n18917 a_43892_n18820 VDD.t2414 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3690 VDD.t1225 a_45772_n17349 a_45684_n17252 VDD.t1224 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3691 a_13623_n12196.t8 a_21772_n14564.t15 VDD.t1878 VDD.t1877 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3692 VDD.t4259 a_26266_n13736 a_26702_n13736 VDD.t4258 pfet_06v0 ad=0.1656p pd=1.28u as=61.199993f ps=0.7u w=0.36u l=0.5u
D106 VSS.t820 a_24481_761.t85 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3693 a_22016_n8961 a_21604_n8548 VSS.t4033 VSS.t4032 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3694 VSS.t2656 a_25544_n16412 a_23564_n11428 VSS.t2655 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X3695 VDD.t1227 a_45772_n14213 a_45684_n14116 VDD.t1226 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3696 VSS.t3076 a_27001_n4328.t2 a_22264_n1148.t0 VSS.t3075 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X3697 VDD.t3594 a_41740_n18917 a_41652_n18820 VDD.t3593 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3698 VDD.t1418 a_43532_n17349 a_43444_n17252 VDD.t1417 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3699 a_28736_n4633.t17 a_30452_n5156.t11 a_31292_n5112 VSS.t1082 nfet_06v0 ad=0.4161p pd=1.905u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3700 VDD.t3820 a_23703_n5156.t7 a_23319_n2759 VDD.t3819 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3701 VDD.t2247 a_23507_n2759 a_25423_n4328 VDD.t2246 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X3702 VDD.t1980 a_40620_n18917 a_40532_n18820 VDD.t1979 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3703 VDD.t1229 a_43532_n14213 a_43444_n14116 VDD.t1228 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3704 VDD.t3080 a_38984_n1975 a_23564_n452.t1 VDD.t3079 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3705 VDD.t196 a_38256_1564.t17 OUT[3].t12 VDD.t195 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3706 a_28744_n14432 a_26532_n14437 a_27804_n14165 VDD.t1959 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X3707 a_43084_n7941 a_42996_n7844 VSS.t2447 VSS.t2446 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3708 a_22052_n4708 a_21604_n5067 VDD.t2066 VDD.t2065 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X3709 a_46220_n6373 a_46132_n6276 VSS.t2086 VSS.t2085 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3710 VDD.t2453 a_26719_n7464 a_27175_n7442 VDD.t2452 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
D107 a_21692_n6694.t23 VDD.t642 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3711 VDD.t1488 a_46556_n1669 a_46468_n1572 VDD.t1158 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3712 a_26999_n10808 a_26543_n11384 VDD.t1949 VDD.t1948 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X3713 VSS.t2576 a_44004_n1192 a_44640_1944.t2 VSS.t2575 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3714 VDD.t770 a_24481_761.t86 a_33467_1116 VDD.t769 pfet_06v0 ad=0.29465p pd=1.74u as=0.26p ps=1.52u w=1u l=0.5u
X3715 a_26440_n5940.t3 a_28156_n6412.t26 VSS.t750 VSS.t749 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3716 a_44092_n7508 a_44004_n7464 VSS.t3275 VSS.t3274 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3717 VSS.t822 a_24481_761.t87 a_30752_1248 VSS.t821 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3718 a_38853_n617 a_38733_n727 VSS.t2024 VSS.t2023 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X3719 a_37484_n15781 a_37396_n15684 VSS.t1375 VSS.t1374 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3720 VSS.t1789 a_37024_1944.t21 OUT[2].t1 VSS.t1788 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3721 VDD.t3611 a_38716_n4805 a_38628_n4708 VDD.t3610 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3722 VSS.t1217 a_23564_n8292 a_21772_n8292.t0 VSS.t1216 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3723 a_26887_n1192 a_26431_n1192 VDD.t3191 VDD.t3190 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X3724 VDD.t3185 a_32650_n12168 a_33086_n12168 VDD.t3184 pfet_06v0 ad=0.1656p pd=1.28u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3725 a_35244_n15781 a_35156_n15684 VSS.t1941 VSS.t1940 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3726 a_23507_n2759 a_22164_n2760 a_23319_n2759 VDD.t1869 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3727 a_24828_n18917 a_24740_n18820 VSS.t3903 VSS.t2637 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3728 a_29161_n14476 a_23072_n13432.t81 VDD.t526 VDD.t525 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X3729 a_37820_n5940 a_37732_n5896 VSS.t1512 VSS.t1511 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3730 a_24684_n16432 a_24964_n14116 a_25559_n10980 VDD.t1836 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3731 VDD.t2846 a_38828_n18917 a_38740_n18820 VDD.t2845 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3732 a_27404_n14990 a_21692_n6694.t24 a_28420_n14820 VSS.t690 nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3733 VDD.t3151 a_28940_n2406.t7 a_29479_n13735 VDD.t3150 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3734 VSS.t4004 a_35064_1506 a_34872_1619 VSS.t4003 nfet_06v0 ad=0.2016p pd=1.48u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3735 a_29612_n8292 a_36773_n5468 a_36709_n5412 VSS.t3170 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3736 VDD.t4301 a_30428_n12645 a_30340_n12548 VDD.t4300 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3737 VDD.t3405 a_34796_n17349 a_34708_n17252 VDD.t3404 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3738 a_34348_n3140 a_34248_n3310 VSS.t2861 VSS.t2860 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3739 a_33832_n8572 a_34092_n9076 VDD.t1775 VDD.t1774 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X3740 VDD.t3315 a_31884_n18917 a_31796_n18820 VDD.t3314 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3741 VDD.t1420 a_34796_n14213 a_34708_n14116 VDD.t1419 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3742 VSS.t1677 a_21772_n452.t13 a_13623_n22908.t6 VSS.t1676 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3743 VSS.t1018 a_26239_n11428 a_26175_n11383 VSS.t1017 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X3744 VDD.t1242 a_32556_n17349 a_32468_n17252 VDD.t1241 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3745 VSS.t1573 a_33077_n1191 a_35940_n1931 VSS.t1572 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3746 a_31628_n5940.t19 a_33496_n6659.t34 VDD.t182 VDD.t181 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3747 a_24771_n2804 a_25547_n2445 a_25139_n2704 VDD.t3892 pfet_06v0 ad=0.1079p pd=0.935u as=0.1826p ps=1.71u w=0.415u l=0.5u
X3748 VSS.t111 a_11023_n6840.t35 a_11087_n7460.t12 VSS.t60 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3749 a_30901_n408 a_30781_n452 VSS.t3400 VSS.t3399 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X3750 VDD.t2171 a_46668_n101 a_46580_n4 VDD.t2170 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3751 VDD.t3680 a_30316_n17349 a_30228_n17252 VDD.t3679 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3752 VDD.t3662 a_23564_n452.t5 a_21772_n452.t0 VDD.t3661 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3753 a_30884_n5112 a_30452_n5156.t12 a_28736_n4633.t16 VSS.t1083 nfet_06v0 ad=0.1312p pd=1.14u as=0.4161p ps=1.905u w=0.82u l=0.6u
X3754 a_37221_n3543 a_36217_n3500 VSS.t1197 VSS.t1196 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X3755 VDD.t3681 a_33900_n15348 a_33812_n15304 VDD.t2385 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3756 a_24693_n9816 a_24573_n9860 a_23949_n9860 VSS.t3943 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X3757 VDD.t1683 a_42748_n10644 a_42660_n10600 VDD.t1682 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3758 a_33533_908 a_24716_1208.t5 VDD.t2187 VDD.t2186 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X3759 a_22772_n4240 a_23072_n13432.t82 VDD.t528 VDD.t527 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X3760 a_21692_n13308.t9 a_26328_n6654.t20 VDD.t2637 VDD.t2636 pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3761 a_29479_n13735 a_30159_n13296 VDD.t3651 VDD.t3650 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3762 VDD.t3454 a_45772_n7941 a_45684_n7844 VDD.t3453 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3763 VDD.t1189 a_43644_n20052 a_43556_n20008 VDD.t1188 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3764 VDD.t1987 a_45772_n4805 a_45684_n4708 VDD.t1986 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3765 VDD.t1801 a_40508_n10644 a_40420_n10600 VDD.t1800 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3766 VSS.t409 a_21692_n5468.t27 a_29444_n708 VSS.t408 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3767 VDD.t950 a_41404_n20052 a_41316_n20008 VDD.t949 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3768 VDD.t3906 a_29408_1944.t21 OUT[0].t10 VDD.t3905 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3769 VSS.t1051 a_21772_n17700.t20 a_13623_n9518.t7 VSS.t1050 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3770 a_42748_n16916 a_42660_n16872 VSS.t1252 VSS.t1251 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3771 a_23072_n13432.t6 a_29744_n15604.t19 VDD.t1645 VDD.t1644 pfet_06v0 ad=0.4392p pd=1.94u as=0.367p ps=1.92u w=1.22u l=0.5u
X3772 a_26440_n5940.t1 a_28156_n6412.t27 VDD.t118 VDD.t117 pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X3773 a_13623_n9518.t5 a_21772_n17700.t21 VSS.t1053 VSS.t1052 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3774 VSS.t1599 a_21772_n14564.t16 a_13623_n12196.t3 VSS.t1598 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3775 VSS.t1256 a_33048_n7420 a_32856_n7376 VSS.t1255 nfet_06v0 ad=0.2016p pd=1.48u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3776 a_30348_n8548 a_29900_n10600.t7 a_29532_n4372.t3 VSS.t3946 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3777 a_25500_n10644 a_25412_n10600 VSS.t2230 VSS.t2229 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3778 a_40508_n16916 a_40420_n16872 VSS.t2712 VSS.t2711 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3779 a_13623_n12196.t2 a_21772_n14564.t17 VSS.t1601 VSS.t1600 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3780 a_36112_n3456 a_34000_n3140 a_35800_n3456 VDD.t2705 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X3781 VDD.t2994 a_27001_n4328.t3 a_22264_n1148.t1 VDD.t2993 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3782 VSS.t1086 a_33494_n9860 a_21916_n6694.t0 VSS.t1085 nfet_06v0 ad=0.2911p pd=1.53u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3783 VDD.t2580 a_41852_n18484 a_41764_n18440 VDD.t2579 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D108 a_25940_n17606.t20 VDD.t4121 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3784 a_31525_n408 a_31405_n452 a_30781_n452 VSS.t3348 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X3785 VDD.t1460 a_33292_n2716 a_33188_n2672 VDD.t1459 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3786 VDD.t2919 a_23564_n3588.t8 a_21772_n3588.t3 VDD.t2918 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3787 a_31968_n704 a_29856_n1121 a_31656_n704 VDD.t943 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X3788 a_33077_n1191 a_32073_n844 VDD.t3018 VDD.t3017 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X3789 VSS.t3767 a_24569_n11820 a_24464_n11680 VSS.t3766 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X3790 a_13623_n4162.t12 a_21772_1116.t15 VDD.t454 VDD.t453 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3791 a_32308_n1976 a_29532_n4372.t7 a_32100_n1976 VSS.t2124 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3792 VSS.t1313 a_21804_n2273.t12 a_21716_n2229 VSS.t1312 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3793 a_10712_4516.t9 a_3935_4156.t14 VSS.t463 VSS.t376 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3794 OUT[4].t1 a_41392_1944.t22 VSS.t1440 VSS.t1439 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3795 VDD.t3463 a_37221_n3543 a_40196_n1884 VDD.t3462 pfet_06v0 ad=0.35315p pd=1.96u as=0.2486p ps=2.01u w=0.565u l=0.5u
X3796 a_30555_n2729 a_29900_n10600.t8 a_30759_n2276 VSS.t3947 nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X3797 VDD.t2075 a_26383_1944 a_26839_1966 VDD.t2074 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X3798 a_29537_n14432 a_23072_n13432.t83 VSS.t534 VSS.t533 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X3799 VDD.t1570 a_24233_n13388 a_24128_n13248 VDD.t1569 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X3800 VSS.t3467 XRST.t3 a_27540_n20747 VSS.t3466 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X3801 a_24609_n3840 a_23072_n13432.t84 VSS.t536 VSS.t535 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X3802 VSS.t538 a_23072_n13432.t85 a_29699_n6600 VSS.t537 nfet_06v0 ad=0.1224p pd=1.04u as=0.134p ps=1.1u w=0.36u l=0.6u
X3803 a_29479_n13735 a_28121_n10980 a_27820_n16432 VDD.t3597 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3804 a_42277_n616 a_42157_n660 a_41533_n727 VSS.t1799 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X3805 a_27001_n4328.t1 a_26271_n4306 VDD.t2852 VDD.t2851 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X3806 VDD.t4071 a_23619_n9860 a_22264_n10556 VDD.t4070 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3807 VDD.t1617 a_46556_n16916 a_46468_n16872 VDD.t1616 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3808 VDD.t152 a_31628_n5940.t42 a_29800_n5940.t3 VDD.t151 pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X3809 a_26635_n12996 a_26983_n12728 VDD.t3888 VDD.t3887 pfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X3810 a_23542_n1754 a_23954_n2020 a_24074_n1976 VSS.t2279 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3811 VSS.t598 a_13623_n4162.t38 a_11023_n4162.t2 VSS.t597 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3812 a_39164_n4372 a_39076_n4328 VSS.t2869 VSS.t2868 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3813 VDD.t1260 a_46556_n13780 a_46468_n13736 VDD.t1259 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3814 VSS.t2045 a_30320_n6636 a_30215_n6265 VSS.t2044 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3815 VDD.t1402 a_32668_n20052 a_32580_n20008 VDD.t1401 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3816 a_45884_n20485 a_45796_n20388 VSS.t2399 VSS.t2398 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3817 a_25139_n2704 a_23072_n13432.t86 a_25159_n2276 VSS.t539 nfet_06v0 ad=0.3123p pd=2.38u as=48.6f ps=0.645u w=0.405u l=0.6u
X3818 a_11087_n10138.t15 a_11023_n9518.t35 a_13501_n9138.t7 VDD.t548 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3819 OUT[5].t5 a_44640_1944.t18 VSS.t270 VSS.t269 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3820 a_35064_1506 a_34576_1204 a_35324_1564 VDD.t1565 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3821 a_41203_n799 a_41533_n727 a_41653_n617 VSS.t3637 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X3822 a_2167_3472.t38 a_11023_n4162.t35 VSS.t2765 VDD.t2698 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3823 a_26981_n10025 a_26861_n10135 VSS.t1619 VSS.t1618 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X3824 VDD.t3442 a_42188_n18917 a_42100_n18820 VDD.t3441 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3825 VDD.t772 a_24481_761.t88 a_29744_n15604.t3 VDD.t771 pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X3826 VDD.t2124 a_42412_n5940 a_42324_n5896 VDD.t2123 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3827 VDD.t1406 a_30428_n20052 a_30340_n20008 VDD.t1405 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3828 a_33496_n6659.t7 CLK.t13 VSS.t2076 VSS.t2075 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X3829 a_42524_n20485 a_42436_n20388 VSS.t2405 VSS.t2404 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3830 VSS.t1369 a_13623_n14874.t39 a_11023_n14874.t15 VSS.t1368 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X3831 OUT[2].t0 a_37024_1944.t22 VSS.t1791 VSS.t1790 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3832 a_29771_n1976 a_29295_n1400 a_29519_n1976 VSS.t1541 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X3833 VDD.t1911 a_38716_n9076 a_38628_n9032 VDD.t1910 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3834 a_46556_n20052 a_46468_n20008 VSS.t3477 VSS.t3476 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3835 a_39357_n660 a_30732_332.t5 VDD.t1604 VDD.t1603 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X3836 a_40508_n7508 a_40420_n7464 VSS.t2780 VSS.t2779 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3837 VDD.t3601 a_25880_n11708 a_21692_n5111.t1 VDD.t3600 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3838 a_11023_n14874.t16 a_13623_n14874.t40 VSS.t1371 VSS.t1370 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3839 VDD.t1469 a_26736_n364 a_26631_7 VDD.t1468 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X3840 a_26747_n1976 a_26271_n1400 a_26495_n1976 VSS.t2581 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X3841 a_29196_n18917 a_29108_n18820 VSS.t2585 VSS.t2584 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3842 a_33029_951 a_32909_841 VSS.t4314 VSS.t4313 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X3843 a_46668_n9509 a_46580_n9412 VSS.t4345 VSS.t4344 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3844 VDD.t2221 a_30876_n18484 a_30788_n18440 VDD.t2220 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3845 VSS.t1901 a_37785_n364 a_37680_n320 VSS.t1900 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X3846 a_24751_n3544 a_24631_n3588 VSS.t3309 VSS.t3308 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X3847 a_21772_n20836.t5 a_23564_n20836 VDD.t885 VDD.t884 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3848 VSS.t96 a_13623_n17552.t37 a_11023_n17552.t2 VSS.t95 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3849 a_42168_1564 a_41616_1564 a_41964_1564 VDD.t2746 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3850 a_11087_n7460.t21 a_11023_n6840.t36 a_13501_n6460.t7 VDD.t115 pfet_03v3 ad=0.728p pd=3.32u as=1.82p ps=6.9u w=2.8u l=0.28u
X3851 VDD.t654 a_21772_n20836.t21 a_13623_n6840.t10 VDD.t653 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3852 a_11087_n23528.t51 a_2167_3472.t51 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X3853 a_11023_n17552.t1 a_13623_n17552.t38 VSS.t98 VSS.t97 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X3854 VDD.t350 a_26388_n17606.t10 a_22220_690.t1 VDD.t349 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3855 a_22052_1944 a_21604_2475 VSS.t2384 VSS.t2383 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
D109 a_23072_n13432.t87 VDD.t529 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3856 a_37372_n18484 a_37284_n18440 VSS.t4019 VSS.t4018 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3857 a_28048_1248 a_25936_1564 a_27736_1248 VDD.t1427 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X3858 a_21692_n13308.t8 a_26328_n6654.t21 VDD.t2639 VDD.t2638 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3859 VSS.t200 a_11023_n22908.t36 a_11087_n23528.t21 VSS.t60 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3860 VSS.t824 a_24481_761.t89 a_26944_1248 VSS.t823 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3861 a_13623_n22908.t7 a_21772_n452.t14 VSS.t1679 VSS.t1678 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3862 VSS.t3097 a_32073_n844 a_31968_n704 VSS.t3096 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X3863 a_42188_n4805 a_42100_n4708 VSS.t1494 VSS.t1493 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3864 a_36252_n18484 a_36164_n18440 VSS.t3936 VSS.t3935 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3865 a_37372_n15348 a_37284_n15304 VSS.t1245 VSS.t1244 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3866 VDD.t2267 a_36140_n13780 a_36052_n13736 VDD.t2266 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3867 a_39164_n13780 a_39076_n13736 VSS.t3835 VSS.t3834 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3868 a_24128_n8544 a_21604_n8548 a_23816_n8544 VSS.t4031 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3869 a_45324_n3237 a_45236_n3140 VSS.t2741 VSS.t2740 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3870 a_39164_n10644 a_39076_n10600 VSS.t2176 VSS.t2175 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3871 a_27643_n11384 a_27167_n10808 a_27391_n11384 VSS.t3657 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X3872 a_45648_1564.t1 a_40652_n1572 VSS.t923 VSS.t922 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3873 a_24128_n5408 a_21604_n5412 a_23816_n5408 VSS.t3579 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3874 VSS.t1845 a_13623_n12196.t40 a_11023_n12196.t16 VSS.t1844 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X3875 a_34012_n18484 a_33924_n18440 VSS.t3932 VSS.t3931 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3876 a_43980_n17349 a_43892_n17252 VSS.t1140 VSS.t1139 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3877 a_26523_n3753 a_26047_n4328 a_26271_n4306 VSS.t2646 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X3878 a_11023_n12196.t17 a_13623_n12196.t41 VSS.t1847 VSS.t1846 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3879 a_11087_n23528.t52 a_2167_3472.t50 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X3880 VDD.t3485 a_33900_n17349 a_33812_n17252 VDD.t3484 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3881 a_43980_n14213 a_43892_n14116 VSS.t953 VSS.t952 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3882 VSS.t1010 a_39056_820 a_38951_420 VSS.t1009 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3883 a_43196_n4372 a_43108_n4328 VSS.t3996 VSS.t3995 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3884 a_22876_n8988 a_22568_n8944 VSS.t3757 VSS.t3756 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X3885 VDD.t2797 a_28524_n18484 a_28436_n18440 VDD.t2796 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3886 a_24731_n3124.t0 a_25019_n3588.t6 VDD.t3392 VDD.t2687 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3887 a_41740_n17349 a_41652_n17252 VSS.t1292 VSS.t1291 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3888 VDD.t4079 a_33900_n14213 a_33812_n14116 VDD.t4078 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3889 VDD.t2714 a_22052_1944 a_29408_1944.t5 VDD.t2713 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3890 a_32108_n2332.t0 a_35456_n4628.t21 VSS.t4171 VSS.t4170 nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X3891 a_22876_n5852 a_22568_n5808 VSS.t1063 VSS.t1062 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X3892 VSS.t2642 a_24573_n12996 a_24693_n12952 VSS.t2641 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3893 a_40620_n17349 a_40532_n17252 VSS.t1296 VSS.t1295 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3894 a_41740_n14213 a_41652_n14116 VSS.t1298 VSS.t1297 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3895 a_11087_n18172.t36 a_2167_3472.t74 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X3896 a_40620_n14213 a_40532_n14116 VSS.t1422 VSS.t1421 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3897 a_24128_n13248 a_22016_n13665 a_23816_n13248 VDD.t3849 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X3898 VDD.t976 a_42748_n9076 a_42660_n9032 VDD.t975 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3899 a_31799_n7508 a_32455_n7420 a_32351_n7376 VDD.t4260 pfet_06v0 ad=0.25375p pd=1.51u as=0.1313p ps=1.025u w=0.505u l=0.5u
D110 VSS.t4194 a_25940_n17606.t21 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3900 a_31548_n20485 a_31460_n20388 VSS.t4327 VSS.t4326 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3901 VDD.t1394 a_36588_n15348 a_36500_n15304 VDD.t988 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3902 VDD.t3298 a_42412_n101 a_42324_n4 VDD.t3297 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3903 a_45212_n4372 a_45124_n4328 VSS.t3921 VSS.t3920 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3904 a_29699_n6600 a_29559_n6456 a_29211_n6724 VSS.t2977 nfet_06v0 ad=0.134p pd=1.1u as=0.176p ps=1.68u w=0.4u l=0.6u
X3905 VDD.t2523 a_48012_n7941 a_47924_n7844 VDD.t2522 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3906 a_23360_n15233 a_22948_n14820 VDD.t2034 VDD.t2033 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X3907 a_27736_1248 a_25936_1564 a_26796_1515 VSS.t1485 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X3908 a_11087_n7460.t11 a_11023_n6840.t37 VSS.t112 VSS.t62 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3909 VDD.t2248 a_34460_n20485 a_34372_n20388 VDD.t2218 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3910 a_2167_3472.t8 a_13623_n4162.t39 VSS.t600 VSS.t599 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X3911 VDD.t2250 a_48012_n4805 a_47924_n4708 VDD.t2249 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3912 VDD.t3183 a_22876_n8988 a_22772_n8944 VDD.t3182 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3913 VSS.t637 a_13623_n20230.t38 a_11023_n20230.t1 VSS.t636 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3914 VDD.t1329 a_34348_n15348 a_34260_n15304 VDD.t1328 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3915 a_27484_n4 a_27032_51 VDD.t865 VDD.t864 pfet_06v0 ad=0.2028p pd=1.3u as=0.45p ps=2.02u w=0.78u l=0.5u
X3916 VDD.t3000 a_22876_n5852 a_22772_n5808 VDD.t2999 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3917 a_47564_n12645 a_47476_n12548 VSS.t4284 VSS.t4283 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3918 a_23072_n13432.t7 a_29744_n15604.t20 VDD.t1647 VDD.t1646 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3919 VDD.t1127 a_25084_1564 a_33216_1944.t6 VDD.t1126 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3920 a_26488_1564 a_25524_1243 a_26284_1564 VSS.t1415 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3921 VSS.t3501 a_43833_1204 a_43728_1248 VSS.t3500 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X3922 a_11023_n22908.t1 a_13623_n22908.t30 VSS.t226 VSS.t225 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3923 a_27496_n14116 a_26532_n14437 a_27292_n14116 VSS.t2034 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X3924 VSS.t2453 a_25795_n2716.t5 a_25547_n2445 VSS.t847 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3925 VDD.t3272 a_31100_n20485 a_31012_n20388 VDD.t3271 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3926 OUT[3].t11 a_38256_1564.t18 VDD.t198 VDD.t197 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3927 a_25940_n17606.t1 a_32262_n452 VDD.t1391 VDD.t1390 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X3928 a_45324_n12645 a_45236_n12548 VSS.t4288 VSS.t4287 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3929 VSS.t228 a_13623_n22908.t31 a_11023_n22908.t0 VSS.t227 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3930 a_40196_1944 a_39748_2475 VSS.t1547 VSS.t1546 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X3931 a_37585_n3140 a_22220_690.t14 a_37605_n3544 VSS.t837 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X3932 VDD.t1665 a_23564_n11428 a_21772_n11428.t4 VDD.t1664 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3933 a_42948_n1976 a_42244_n1572 VSS.t3877 VSS.t3876 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3934 a_34708_n5896.t8 a_33776_n5896.t20 VDD.t842 VDD.t841 pfet_06v0 ad=0.4392p pd=1.94u as=0.367p ps=1.92u w=1.22u l=0.5u
X3935 a_25276_n18484 a_25188_n18440 VSS.t3630 VSS.t3629 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D111 VSS.t540 a_23072_n13432.t88 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3936 a_13623_n14874.t11 a_21772_n11428.t20 VDD.t310 VDD.t309 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3937 a_24388_n4708 a_21916_n6694.t18 VDD.t1065 VDD.t1064 pfet_06v0 ad=0.3782p pd=1.84u as=0.6588p ps=3.52u w=1.22u l=0.5u
X3938 VDD.t2897 a_46668_n11077 a_46580_n10980 VDD.t2896 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3939 a_11087_n23528.t53 a_2167_3472.t49 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X3940 a_38828_n17349 a_38740_n17252 VSS.t3458 VSS.t3457 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3941 a_33188_n2672 a_24481_761.t90 VDD.t774 VDD.t773 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X3942 VDD.t312 a_21772_n11428.t21 a_13623_n14874.t10 VDD.t311 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3943 a_23036_n18484 a_22948_n18440 VSS.t3656 VSS.t3655 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3944 a_38828_n14213 a_38740_n14116 VSS.t3463 VSS.t3462 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3945 VDD.t1631 a_42860_n5940 a_42772_n5896 VDD.t1630 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3946 a_11087_n10138.t28 a_13623_n9518.t31 a_13501_n9138.t11 VSS.t263 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3947 a_25836_n1236.t5 a_34649_n2412 VDD.t3621 VDD.t3620 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3948 VDD.t3199 a_44428_n11077 a_44340_n10980 VDD.t3198 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3949 VDD.t4241 a_26563_n12212 a_26431_n12168 VDD.t4240 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X3950 VSS.t2689 a_21692_n13308.t30 a_22948_n14820 VSS.t2688 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X3951 a_40060_n4805 a_39972_n4708 VSS.t1995 VSS.t1994 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3952 a_33784_n6976 a_32856_n7376 a_33616_n6976 VSS.t2826 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3953 a_25880_n11708 a_25860_n9032 VDD.t2077 VDD.t2076 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X3954 VSS.t1656 a_32413_n14564 a_32533_n14520 VSS.t1655 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3955 a_40956_n7508 a_40868_n7464 VSS.t4256 VSS.t4255 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3956 a_11087_n23528.t54 a_2167_3472.t48 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X3957 a_30764_n17349 a_30676_n17252 VSS.t3465 VSS.t3464 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D112 VSS.t541 a_23072_n13432.t89 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X3958 VSS.t3792 a_25132_n16432 a_23608_n15260 VSS.t3791 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X3959 a_11087_n20850.t22 a_13623_n20230.t39 a_13501_n19850.t12 VSS.t638 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3960 VDD.t322 a_26440_n5940.t16 a_21692_n5468.t8 VDD.t321 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X3961 a_13623_n22908.t0 a_21772_n452.t15 VDD.t1598 VDD.t1597 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3962 a_22568_n8944 a_22016_n8961 a_22364_n8944 VDD.t3785 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3963 a_30752_n11296 a_30604_n11029 a_30584_n11296 VSS.t1518 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3964 a_48012_n15781 a_47924_n15684 VSS.t2082 VSS.t2081 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3965 VSS.t272 a_44640_1944.t19 OUT[5].t4 VSS.t271 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3966 a_23038_n1422 a_22918_n2020 VDD.t4037 VDD.t4036 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X3967 a_43868_n1669 a_43780_n1572 VSS.t3380 VSS.t2400 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3968 a_36520_n3868 a_10712_4516.t49 VSS.t353 VSS.t352 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X3969 a_28617_n8548 a_24492_n5156 a_28433_n8548 VSS.t3584 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X3970 a_13501_n22528.t2 a_13623_n22908.t32 a_11087_n23528.t2 VSS.t229 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X3971 VDD.t3424 a_47900_n16916 a_47812_n16872 VDD.t3423 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3972 a_22568_n5808 a_22016_n5825 a_22364_n5808 VDD.t3072 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3973 a_41852_n12212 a_41764_n12168 VSS.t3711 VSS.t3710 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3974 a_11087_n23528.t55 a_2167_3472.t47 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X3975 VDD.t2785 a_36428_n53 a_36324_n4 VDD.t2784 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3976 a_21772_n17700.t4 a_23564_n17700 VDD.t4243 VDD.t4242 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3977 VDD.t1740 a_47900_n13780 a_47812_n13736 VDD.t1739 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3978 VDD.t2822 a_45772_n18917 a_45684_n18820 VDD.t2821 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3979 VDD.t3806 a_47564_n17349 a_47476_n17252 VDD.t3805 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3980 VDD.t4004 a_29308_n20485 a_29220_n20388 VDD.t4003 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3981 a_21772_n14564.t2 a_23564_n14564.t7 VDD.t3744 VDD.t3743 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X3982 VSS.t1681 a_21772_n452.t16 a_13623_n22908.t5 VSS.t1680 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3983 a_39408_n4 a_39308_n452 VDD.t2672 VDD.t2671 pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X3984 a_23024_n3840 a_22876_n4284 a_22856_n3840 VSS.t3410 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3985 VSS.t2946 a_27597_n8292 a_27717_n8248 VSS.t2945 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X3986 VDD.t3470 a_47564_n14213 a_47476_n14116 VDD.t3469 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3987 a_45772_n3237 a_45684_n3140 VSS.t1665 VSS.t1664 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3988 a_27988_n4328 a_27540_n3797 VDD.t2181 VDD.t2180 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X3989 VDD.t3105 a_23703_n5156.t8 a_23207_n4708 VDD.t3104 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X3990 VDD.t822 a_34708_n5896.t27 a_35456_n4628.t4 VDD.t821 pfet_06v0 ad=0.367p pd=1.92u as=0.2952p ps=1.54u w=0.82u l=0.5u
X3991 VDD.t3713 a_43532_n18917 a_43444_n18820 VDD.t3712 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D113 a_23072_n13432.t90 VDD.t530 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X3992 a_23016_n7376 a_22464_n7393 a_22812_n7376 VDD.t4045 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X3993 a_33832_n8572 a_34092_n9076 VSS.t1861 VSS.t1860 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X3994 VDD.t3111 a_45324_n17349 a_45236_n17252 VDD.t3110 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3995 VDD.t3113 a_45324_n14213 a_45236_n14116 VDD.t3112 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X3996 VSS.t186 a_38256_1564.t19 OUT[3].t1 VSS.t185 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X3997 a_47900_n20052 a_47812_n20008 VSS.t3889 VSS.t3888 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X3998 a_11087_n10138.t30 a_2167_3472.t83 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X3999 a_37932_n9509 a_37844_n9412 VSS.t3469 VSS.t3468 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4000 a_35468_n12645 a_35380_n12548 VSS.t1538 VSS.t1537 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4001 VDD.t3478 a_38380_n15781 a_38292_n15684 VDD.t3477 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4002 a_25836_n1236.t4 a_34649_n2412 VDD.t3619 VDD.t3618 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X4003 a_11023_n4162.t1 a_13623_n4162.t40 VSS.t602 VSS.t601 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4004 a_27804_n14165 a_27496_n14116 VSS.t2052 VSS.t2051 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X4005 VDD.t3685 a_37260_n12645 a_37172_n12548 VDD.t3684 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4006 VDD.t4050 a_36140_n15781 a_36052_n15684 VDD.t2776 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4007 a_28300_n18917 a_28212_n18820 VSS.t3000 VSS.t2999 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4008 VSS.t35 a_45648_1564.t18 EOC.t4 VSS.t34 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4009 VSS.t705 a_29800_n5940.t20 a_28156_n6412.t2 VSS.t704 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X4010 VDD.t3294 a_42972_n1236 a_42884_n1192 VDD.t3293 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4011 VDD.t3016 a_35020_n12645 a_34932_n12548 VDD.t3015 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D114 a_21692_n6694.t25 VDD.t643 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X4012 VDD.t3908 a_29408_1944.t22 OUT[0].t9 VDD.t3907 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4013 a_27225_n1572.t0 a_26495_n1976 VSS.t2481 VSS.t2480 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X4014 a_45660_n4372 a_45572_n4328 VSS.t3998 VSS.t3997 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4015 VDD.t1606 a_30732_332.t6 a_30576_376 VDD.t1605 pfet_06v0 ad=0.4392p pd=1.94u as=0.4758p ps=2u w=1.22u l=0.5u
X4016 VSS.t1104 a_21916_n6694.t19 a_21812_n6643 VSS.t1103 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X4017 a_39276_n15781 a_39188_n15684 VSS.t4242 VSS.t4241 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4018 VDD.t4067 a_37260_n7941 a_37172_n7844 VDD.t4066 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4019 VSS.t3829 a_29540_n11728 a_24492_n5156 VSS.t3828 nfet_06v0 ad=0.224p pd=1.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4020 a_37036_n15781 a_36948_n15684 VSS.t3729 VSS.t3728 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4021 VDD.t1923 a_46108_n7508 a_46020_n7464 VDD.t1922 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4022 a_32309_n9240 a_32189_n9860 a_31565_n9860 VDD.t2654 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X4023 VSS.t2747 a_24403_n2414 a_24315_n2759 VSS.t2746 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X4024 VDD.t2357 a_25795_n2716.t6 a_25547_n2445 VDD.t2356 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X4025 VDD.t3822 a_46108_n4372 a_46020_n4328 VDD.t3821 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4026 VDD.t3672 a_35804_n16916 a_35716_n16872 VDD.t3671 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4027 a_35568_n4 a_35156_n325 VDD.t2985 VDD.t2984 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X4028 VDD.t3878 a_34796_n18917 a_34708_n18820 VDD.t3877 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4029 VDD.t2534 a_36588_n17349 a_36500_n17252 VDD.t2533 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4030 a_26271_n1400 a_25647_n1976 a_26123_n1976 VSS.t1996 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4031 a_21996_n12996.t0 a_30584_n1954 VSS.t3598 VSS.t3597 nfet_06v0 ad=0.1261p pd=1.005u as=0.2134p ps=1.85u w=0.485u l=0.6u
X4032 a_23479_n5156 a_26943_n7442 VDD.t2887 VDD.t2886 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X4033 a_41516_n5940 a_41428_n5896 VSS.t1704 VSS.t1703 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4034 VDD.t4137 a_36588_n14213 a_36500_n14116 VDD.t2323 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4035 VDD.t2538 a_34348_n17349 a_34260_n17252 VDD.t2537 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4036 a_28972_n7819 a_28852_n8292.t3 VDD.t3581 VDD.t3580 pfet_06v0 ad=0.2847p pd=1.615u as=0.5913p ps=3.27u w=1.095u l=0.5u
X4037 a_25795_n2716.t0 a_21692_n5468.t28 VSS.t371 VSS.t370 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4038 a_22772_n4240 a_21604_n3844 a_22568_n4240 VDD.t1714 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X4039 VDD.t3181 a_31436_n18917 a_31348_n18820 VDD.t3180 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4040 a_42188_n17349 a_42100_n17252 VSS.t1001 VSS.t1000 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4041 VDD.t4140 a_34348_n14213 a_34260_n14116 VDD.t4139 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4042 a_24609_n704 a_23072_n13432.t91 VSS.t543 VSS.t542 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X4043 VDD.t3810 a_32108_n17349 a_32020_n17252 VDD.t3809 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4044 a_42188_n14213 a_42100_n14116 VSS.t1003 VSS.t1002 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4045 VSS.t3317 a_24731_n3124.t4 a_37499_860 VSS.t3316 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X4046 VSS.t2636 a_41203_n799 a_39308_n452 VSS.t2635 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4047 a_35804_n20052 a_35716_n20008 VSS.t3564 VSS.t3563 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4048 VSS.t1450 a_34895_n1192 a_35371_n617 VSS.t1449 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X4049 a_31548_n10172.t9 a_33496_n8222.t20 VDD.t298 VDD.t297 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4050 VDD.t3541 a_24233_n844 a_24128_n704 VDD.t3540 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X4051 VSS.t170 a_33496_n6659.t35 a_31628_n5940.t1 VSS.t169 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X4052 a_29980_n18484 a_29892_n18440 VSS.t2347 VSS.t2346 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4053 a_22016_n13665 a_21604_n13252 VDD.t2139 VDD.t2138 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X4054 VDD.t3397 a_46556_n20052 a_46468_n20008 VDD.t3396 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4055 VDD.t231 a_13623_n22908.t33 a_11023_n22908.t12 VDD.t230 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4056 VSS.t334 a_26440_n5940.t17 a_21692_n5468.t2 VSS.t333 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X4057 a_22016_n10529 a_21604_n10116 VDD.t3365 VDD.t3364 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X4058 OUT[5].t3 a_44640_1944.t20 VSS.t274 VSS.t273 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4059 a_29076_n8292.t0 a_24815_n3588.t18 VDD.t36 VDD.t35 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4060 VDD.t3812 a_41292_n7941 a_41204_n7844 VDD.t3811 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4061 a_30808_n10600 a_29076_n8292.t9 a_30808_n10116 VDD.t441 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4062 a_32413_n12996 a_28927_n10160 VDD.t2310 VDD.t2309 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X4063 VDD.t3209 a_24380_n18917 a_24292_n18820 VDD.t1607 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4064 VSS.t2372 a_30192_n15304.t18 a_24481_761.t6 VSS.t2371 nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X4065 a_38847_464 a_37947_332 VDD.t3282 VDD.t3281 pfet_06v0 ad=0.1313p pd=1.025u as=0.29465p ps=1.74u w=0.505u l=0.5u
X4066 VDD.t2559 a_41292_n4805 a_41204_n4708 VDD.t2558 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4067 VSS.t4060 a_29532_n10311 a_29444_n10116 VSS.t4059 nfet_06v0 ad=0.2344p pd=1.56u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4068 a_26328_n6654.t3 a_28156_n6412.t28 VDD.t120 VDD.t119 pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X4069 a_31235_n9860 a_31565_n9860 a_31685_n9816 VSS.t2290 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
D115 VSS.t691 a_21692_n6694.t26 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X4070 a_24481_761.t4 a_30192_n15304.t19 VSS.t2374 VSS.t2373 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X4071 a_31636_n2760 a_25019_n3588.t7 a_31392_n2760 VDD.t3393 pfet_06v0 ad=0.3172p pd=1.74u as=0.4248p ps=1.94u w=1.22u l=0.5u
X4072 a_21772_n17700.t1 a_23564_n17700 VSS.t4308 VSS.t4307 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4073 VDD.t2114 a_22140_n18917 a_22052_n18820 VDD.t1609 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4074 VSS.t1055 a_21772_n17700.t22 a_13623_n9518.t1 VSS.t1054 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4075 a_21772_n14564.t3 a_23564_n14564.t8 VSS.t3814 VSS.t3813 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4076 a_22364_n4240 a_21792_n7464 VDD.t1028 VDD.t1027 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X4077 VDD.t919 a_43644_n18484 a_43556_n18440 VDD.t918 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4078 VSS.t1603 a_21772_n14564.t18 a_13623_n12196.t1 VSS.t1602 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4079 VSS.t4291 a_43555_n452 a_41864_1394 VSS.t4290 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4080 a_28583_n3140 a_29263_n3588.t3 VDD.t3235 VDD.t3234 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4081 VDD.t2547 a_40172_n9509 a_40084_n9412 VDD.t2546 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4082 a_38256_1564.t4 a_37844_1564 VDD.t4186 VDD.t4185 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4083 VSS.t4260 a_37844_1564 a_38256_1564.t0 VSS.t4259 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4084 VDD.t2553 a_41740_n6373 a_41652_n6276 VDD.t2552 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4085 VDD.t3918 a_41404_n18484 a_41316_n18440 VDD.t3917 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4086 a_22568_n13648 a_22016_n13665 a_22364_n13648 VDD.t3848 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X4087 a_21772_n452.t2 a_23564_n452.t6 VSS.t3745 VSS.t3744 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4088 a_25975_n184 a_26631_7 a_26527_51 VDD.t1429 pfet_06v0 ad=0.25375p pd=1.51u as=0.1313p ps=1.025u w=0.505u l=0.5u
X4089 VDD.t3086 a_41740_n3237 a_41652_n3140 VDD.t3085 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4090 VDD.t1623 a_30555_n13780 a_28927_n10160 VDD.t1622 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X4091 VSS.t3737 a_30159_n13296 a_30095_n13252 VSS.t3736 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X4092 a_27496_n14116 a_26944_n14116 a_27292_n14116 VDD.t3920 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X4093 a_46108_n1669 a_46020_n1572 VSS.t2278 VSS.t1270 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4094 VDD.t2836 a_37372_n12212 a_37284_n12168 VDD.t2835 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D116 VSS.t544 a_23072_n13432.t92 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X4095 VSS.t546 a_23072_n13432.t93 a_30864_n704 VSS.t545 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4096 VDD.t3370 a_36252_n12212 a_36164_n12168 VDD.t3369 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4097 VDD.t592 a_13623_n20230.t40 a_11023_n20230.t12 VDD.t591 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4098 a_38853_n5874 a_38733_n5431 VDD.t2164 VDD.t2163 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X4099 a_35392_n10172 a_34652_n11391 VSS.t4224 VSS.t4223 nfet_06v0 ad=0.1584p pd=1.6u as=0.2344p ps=1.56u w=0.36u l=0.6u
X4100 a_30752_1248 a_30604_1515 a_30584_1248 VSS.t962 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4101 a_44509_n452 a_42948_n1976 VDD.t2988 VDD.t2987 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X4102 a_24828_n20052 a_24740_n20008 VSS.t2638 VSS.t2637 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4103 a_13501_n19850.t1 a_11023_n20230.t36 a_11087_n20850.t16 VDD.t1904 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4104 VDD.t2712 a_22052_1944 a_29408_1944.t4 VDD.t2711 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4105 a_38853_n2738 a_38733_n2295 VDD.t2749 VDD.t2748 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X4106 a_48012_n3237 a_47924_n3140 VSS.t4358 VSS.t4357 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4107 a_28156_n6412.t1 a_29800_n5940.t21 VSS.t707 VSS.t706 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X4108 a_36812_n12645 a_36724_n12548 VSS.t3539 VSS.t3538 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4109 VDD.t1913 a_46556_n7508 a_46468_n7464 VDD.t1912 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4110 a_38604_n7941 a_38516_n7844 VSS.t1137 VSS.t1136 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4111 a_47676_n20485 a_47588_n20388 VSS.t3781 VSS.t3780 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4112 a_11023_n9518.t1 a_13623_n9518.t32 VSS.t265 VSS.t264 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4113 VDD.t3996 a_46108_n16916 a_46020_n16872 VDD.t3995 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4114 a_22588_n2020 a_22918_n2020 a_23038_n1422 VDD.t4035 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X4115 VDD.t2364 a_46556_n4372 a_46468_n4328 VDD.t2363 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4116 VDD.t2561 a_46108_n13780 a_46020_n13736 VDD.t2560 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4117 VDD.t448 a_21772_1116.t16 a_13623_n4162.t11 VDD.t447 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4118 a_45436_n20485 a_45348_n20388 VSS.t3577 VSS.t3576 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4119 VSS.t1321 a_33252_n1192 a_29900_760.t0 VSS.t1320 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4120 a_41964_n5940 a_41876_n5896 VSS.t2701 VSS.t2700 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4121 a_39357_n5364 a_25020_n8200.t6 VDD.t847 VDD.t846 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X4122 a_31405_n452 a_22672_n2214.t4 VSS.t1504 VSS.t1503 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4123 a_31392_n2760 a_31292_n2804 VDD.t2905 VDD.t2904 pfet_06v0 ad=0.4248p pd=1.94u as=0.4972p ps=3.14u w=1.13u l=0.5u
X4124 a_39612_n7508 a_39524_n7464 VSS.t4234 VSS.t4233 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4125 a_39357_n2228 a_37221_n3543 VDD.t3461 VDD.t3460 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X4126 VDD.t3533 a_45212_n1236 a_45124_n1192 VDD.t2548 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4127 VDD.t2629 a_21692_n13308.t31 a_21604_n13252 VDD.t2628 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X4128 VDD.t2631 a_21692_n13308.t32 a_21604_n10116 VDD.t2630 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X4129 a_41616_1564 a_41204_1243 VSS.t1869 VSS.t1868 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4130 a_37368_n320 a_35156_n325 a_36428_n53 VDD.t2983 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X4131 a_46108_n20052 a_46020_n20008 VSS.t2652 VSS.t2651 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4132 VDD.t2272 a_32668_n18484 a_32580_n18440 VDD.t2271 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4133 VDD.t16 a_22444_332.t30 a_27852_n14990 VDD.t15 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X4134 a_13623_n17552.t0 a_21772_n8292.t22 VSS.t47 VSS.t46 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4135 a_27820_n16432 a_28121_n10980 a_29687_n13252 VSS.t3684 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X4136 a_33019_n8457 a_32543_n9032 a_32767_n9010 VSS.t3609 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X4137 a_43644_n705 a_43833_1204 VSS.t3499 VSS.t3498 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X4138 VSS.t4209 a_32108_n2332.t26 a_32020_n2276 VSS.t4208 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X4139 a_42188_n9509 a_42100_n9412 VSS.t1468 VSS.t1467 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4140 a_32880_n10112 a_32732_n10556 a_32712_n10112 VSS.t2154 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4141 VDD.t883 a_23564_n20836 a_21772_n20836.t4 VDD.t882 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4142 VDD.t2274 a_30428_n18484 a_30340_n18440 VDD.t2273 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4143 a_39164_n18484 a_39076_n18440 VSS.t4217 VSS.t4216 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4144 a_34895_376 a_34271_376 a_34727_376 VDD.t3446 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X4145 a_29736_n8548 a_21692_n6694.t27 VSS.t693 VSS.t692 nfet_06v0 ad=0.1722p pd=1.24u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4146 VSS.t3433 a_31459_n12996 a_31279_n11728 VSS.t3432 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4147 VDD.t1649 a_29744_n15604.t21 a_23072_n13432.t7 VDD.t1648 pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X4148 VSS.t363 a_26440_n5940.t18 a_21692_n5468.t1 VSS.t362 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X4149 a_13623_n6840.t9 a_21772_n20836.t22 VDD.t656 VDD.t655 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4150 a_39164_n15348 a_39076_n15304 VSS.t3794 VSS.t3793 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4151 a_38312_n1975 a_22276_n1572.t3 VSS.t4236 VSS.t4235 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X4152 a_38268_n4805 a_38180_n4708 VSS.t4109 VSS.t4108 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4153 VDD.t658 a_21772_n20836.t23 a_13623_n6840.t8 VDD.t657 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4154 VDD.t3139 a_25817_804 a_25137_864 VDD.t3138 pfet_06v0 ad=0.3276p pd=1.62u as=0.2028p ps=1.3u w=0.78u l=0.5u
X4155 a_29360_n12864 a_27744_n12908 a_28232_n12606 VSS.t1568 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4156 VDD.t2604 a_37932_n17349 a_37844_n17252 VDD.t2603 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4157 VDD.t3872 a_38403_n799 a_33820_n452.t1 VDD.t3871 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4158 a_35288_n1975 a_32308_n1976 VSS.t3693 VSS.t3692 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X4159 a_45772_n17349 a_45684_n17252 VSS.t1279 VSS.t1278 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4160 VDD.t2641 a_37932_n14213 a_37844_n14116 VDD.t2640 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4161 a_32189_n9860 a_32581_n9860 VDD.t2842 VDD.t2841 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X4162 VDD.t3172 a_33900_n18917 a_33812_n18820 VDD.t3171 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4163 a_45772_n14213 a_45684_n14116 VSS.t3048 VSS.t3047 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4164 VSS.t2743 a_29161_n14476 a_29056_n14432 VSS.t2742 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X4165 a_42636_n7941 a_42548_n7844 VSS.t4179 VSS.t4178 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4166 a_43532_n17349 a_43444_n17252 VSS.t1474 VSS.t1473 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4167 a_22364_n13648 a_22264_n13692 VDD.t1534 VDD.t1533 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X4168 VDD.t1108 a_21916_n1975 a_21828_n1931 VDD.t1107 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X4169 VDD.t3730 a_25836_n1236.t37 a_22444_332.t0 VDD.t3729 pfet_06v0 ad=0.30535p pd=1.605u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4170 a_25986_n4536 a_25530_n5112 VDD.t3762 VDD.t3761 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X4171 a_25880_n11708 a_25860_n9032 VSS.t2151 VSS.t2150 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X4172 a_43532_n14213 a_43444_n14116 VSS.t3522 VSS.t3521 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4173 VSS.t276 a_44640_1944.t21 OUT[5].t2 VSS.t275 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4174 a_26047_n4328 a_25423_n4328 a_25899_n3752 VSS.t1389 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4175 VDD.t3502 a_27709_n16132 a_27829_n15512 VDD.t3501 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X4176 VDD.t3589 a_27852_n14990 a_26563_n12212 VDD.t3588 pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X4177 a_27292_n14116 a_27192_n14286 VDD.t2467 VDD.t2466 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X4178 a_43644_n7508 a_43556_n7464 VSS.t2072 VSS.t2071 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4179 VDD.t2680 a_42524_n2804 a_42436_n2760 VDD.t2679 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4180 a_38380_n11077 a_38292_n10980 VSS.t2778 VSS.t2777 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4181 a_28736_n4633.t18 a_25836_n1236.t38 VDD.t3732 VDD.t3731 pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X4182 VDD.t3808 a_47900_n20052 a_47812_n20008 VDD.t3807 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4183 VSS.t3368 a_37947_332 a_37859_377 VSS.t3367 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X4184 VDD.t4142 a_22892_n5156.t4 a_22788_n4708 VDD.t4141 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
D117 VSS.t694 a_21692_n6694.t28 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X4185 VDD.t3292 a_37372_n20485 a_37284_n20388 VDD.t2778 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4186 VSS.t1857 a_32579_769 a_28492_332 VSS.t1856 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4187 a_46556_n1669 a_46468_n1572 VSS.t1552 VSS.t1265 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4188 VDD.t3036 a_36252_n20485 a_36164_n20388 VDD.t2094 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4189 a_26839_1966 a_26383_1944 a_26607_1966 VDD.t2073 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X4190 OUT[3].t10 a_38256_1564.t20 VDD.t200 VDD.t199 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4191 VDD.t4023 a_22968_n6679 a_22668_n14864.t1 VDD.t4022 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4192 a_29888_n7464 a_25612_n6679 VDD.t1221 VDD.t1220 pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4193 VDD.t3071 a_41404_n7508 a_41316_n7464 VDD.t3070 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4194 a_11087_n20850.t17 a_11023_n20230.t37 VSS.t1978 VSS.t56 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4195 OUT[3].t0 a_38256_1564.t21 VSS.t188 VSS.t187 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4196 VDD.t1117 a_41404_n4372 a_41316_n4328 VDD.t1116 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4197 VDD.t2856 a_34012_n20485 a_33924_n20388 VDD.t2792 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4198 VDD.t2684 a_29161_n14476 a_29056_n14432 VDD.t2683 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X4199 VSS.t1303 a_33497_n9032 a_34176_n6976 VSS.t1302 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4200 VDD.t2290 a_30192_n15304.t20 a_24481_761.t3 VDD.t1638 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X4201 VSS.t3199 a_28752_n15348 a_27404_n14990 VSS.t3198 nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
X4202 VSS.t3747 a_23564_n452.t7 a_21772_n452.t3 VSS.t3746 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4203 a_47116_n12645 a_47028_n12548 VSS.t3509 VSS.t3508 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4204 a_27709_n16132 a_24348_n16087.t7 VSS.t2516 VSS.t2515 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4205 VSS.t100 a_13623_n17552.t39 a_11023_n17552.t0 VSS.t99 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4206 a_13623_n20230.t9 a_21772_n3588.t16 VDD.t851 VDD.t850 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4207 VDD.t810 a_27259_804.t15 a_22444_332.t1 VDD.t809 pfet_06v0 ad=0.2561p pd=1.505u as=0.52205p ps=2.045u w=0.985u l=0.5u
X4208 a_41292_n12645 a_41204_n12548 VSS.t2166 VSS.t2165 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4209 a_11087_n23528.t20 a_11023_n22908.t37 VSS.t201 VSS.t62 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4210 a_10778_2852.t7 a_10712_4516.t50 VDD.t344 VDD.t343 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4211 a_37024_1944.t4 a_36388_1944 VDD.t1653 VDD.t1652 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4212 a_34367_1619 a_33467_1116 VSS.t3733 VSS.t3732 nfet_06v0 ad=94.5f pd=0.885u as=0.1224p ps=1.04u w=0.36u l=0.6u
X4213 a_31392_n2760 a_25019_n3588.t8 a_31412_n2276 VSS.t3475 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4214 VSS.t2766 a_11023_n4162.t36 VSS.t2766 VSS.t72 nfet_03v3 ad=1.708p pd=6.82u as=0 ps=0 w=2.8u l=0.28u
X4215 a_13623_n4162.t10 a_21772_1116.t17 VDD.t450 VDD.t449 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
D118 VSS.t13 a_22444_332.t31 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X4216 a_41653_n617 a_41533_n727 VSS.t3636 VSS.t3635 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X4217 a_34796_n17349 a_34708_n17252 VSS.t3489 VSS.t3488 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4218 a_36428_n53 a_36120_n4 VDD.t2982 VDD.t2981 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X4219 VSS.t548 a_23072_n13432.t94 a_23472_n6976 VSS.t547 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4220 a_34796_n14213 a_34708_n14116 VSS.t1476 VSS.t1475 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4221 a_41392_1944.t0 a_40196_1944 VSS.t3131 VSS.t3130 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4222 a_2167_3472.t39 a_11023_n4162.t37 VSS.t2767 VDD.t2699 pfet_03v3 ad=1.82p pd=6.9u as=0.728p ps=3.32u w=2.8u l=0.28u
X4223 VSS.t4196 a_25940_n17606.t22 a_26971_n14820 VSS.t4195 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X4224 a_24069_n9262 a_23949_n9860 VDD.t1932 VDD.t1931 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X4225 a_32556_n17349 a_32468_n17252 VSS.t1478 VSS.t1477 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4226 a_30500_1564 a_29332_1243 a_30296_1564 VDD.t2512 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X4227 a_23728_464 a_22724_860.t6 a_23524_464 VSS.t918 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4228 VDD.t3656 a_45660_n1236 a_45572_n1192 VDD.t3037 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4229 a_24152_n11680 a_22352_n12097 a_23212_n12124 VSS.t0 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X4230 a_24069_n6126 a_23949_n6724 VDD.t922 VDD.t921 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X4231 a_11087_n18172.t37 a_2167_3472.t73 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X4232 a_11087_n15494.t8 a_13623_n14874.t41 a_13501_n14494.t8 VSS.t1372 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4233 VDD.t2804 a_36744_n1954 a_30452_n5156.t2 VDD.t2803 pfet_06v0 ad=0.458p pd=2.02u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4234 a_11023_n4162.t0 a_13623_n4162.t41 VSS.t604 VSS.t603 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4235 a_30316_n17349 a_30228_n17252 VSS.t3763 VSS.t3762 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4236 a_33216_1944.t5 a_25084_1564 VDD.t1125 VDD.t1124 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4237 a_34350_n10980 a_22140_n6694.t15 VSS.t4141 VSS.t4140 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X4238 VDD.t3407 a_37820_n7508 a_37732_n7464 VDD.t3406 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4239 a_43644_n12212 a_43556_n12168 VSS.t2909 VSS.t2908 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4240 VDD.t2460 a_27302_n13160 a_27758_n13714 VDD.t2459 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X4241 a_31669_860 a_24631_n3588 VSS.t3307 VSS.t3306 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4242 VDD.t4134 a_32108_n2332.t27 a_32020_n2276 VDD.t4133 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X4243 a_11087_n23528.t56 a_2167_3472.t46 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X4244 VDD.t1346 a_47564_n18917 a_47476_n18820 VDD.t1345 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4245 a_11087_n18172.t2 a_13623_n17552.t40 a_13501_n17172.t2 VSS.t101 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4246 a_30612_n1104 a_23072_n13432.t95 VDD.t532 VDD.t531 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X4247 VDD.t3767 a_21692_2431 a_28671_n1976 VDD.t3766 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X4248 VDD.t3383 a_35804_n20052 a_35716_n20008 VDD.t1002 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4249 VDD.t4279 a_26396_n20485 a_26308_n20388 VDD.t4278 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4250 a_31525_168 a_31405_n452 a_30781_n452 VDD.t3259 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X4251 VDD.t3401 a_47564_n101 a_47476_n4 VDD.t3400 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4252 a_38984_n1975 a_23999_n2320.t6 VDD.t2411 VDD.t2410 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X4253 a_41404_n12212 a_41316_n12168 VSS.t3327 VSS.t3326 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4254 a_26383_n2968 a_25759_n3544 a_26215_n2968 VDD.t3481 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X4255 a_44640_1944.t1 a_44004_n1192 VSS.t2574 VSS.t2573 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4256 VDD.t1322 a_45324_n18917 a_45236_n18820 VDD.t1321 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4257 VDD.t3643 a_47116_n17349 a_47028_n17252 VDD.t3642 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4258 VSS.t743 a_13623_n6840.t40 a_11023_n6840.t17 VSS.t742 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4259 VDD.t3804 a_47900_n9076 a_47812_n9032 VDD.t3803 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4260 a_25767_n11383 a_24964_n14116 VSS.t1909 VSS.t1908 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X4261 a_34908_n16916 a_34820_n16872 VSS.t3520 VSS.t3519 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4262 a_31628_n5940.t0 a_33496_n6659.t36 VSS.t172 VSS.t171 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X4263 VDD.t2064 a_41292_n17349 a_41204_n17252 VDD.t2063 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4264 VDD.t2158 a_47116_n14213 a_47028_n14116 VDD.t2157 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4265 VDD.t2921 a_23564_n3588.t9 a_21772_n3588.t1 VDD.t2920 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4266 a_41292_n3237 a_41204_n3140 VSS.t4066 VSS.t4065 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4267 a_44204_n5940 a_44116_n5896 VSS.t4047 VSS.t4046 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4268 VDD.t2208 a_40172_n17349 a_40084_n17252 VDD.t2207 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4269 VDD.t2173 a_41292_n14213 a_41204_n14116 VDD.t2172 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4270 a_26215_1944 a_25759_1944 VDD.t891 VDD.t890 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X4271 a_11087_n12816.t28 a_13623_n12196.t42 a_13501_n11816.t18 VSS.t1848 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4272 VDD.t357 a_21692_n5468.t29 a_29332_1243 VDD.t356 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X4273 a_28132_376 a_27572_860 a_28004_860 VSS.t1862 nfet_06v0 ad=0.2132p pd=1.34u as=0.1968p ps=1.3u w=0.82u l=0.6u
X4274 VSS.t1575 a_27988_n4328 a_31348_n1931 VSS.t1574 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4275 VDD.t4285 a_30472_n9815 a_25724_n14564 VDD.t4284 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4276 VDD.t1196 a_40172_n14213 a_40084_n14116 VDD.t1195 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4277 a_30092_1564 a_28836_376 VSS.t1697 VSS.t1696 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4278 VDD.t18 a_22444_332.t32 a_27572_860 VDD.t17 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4279 a_40672_864 a_39056_820 a_39544_420 VSS.t1008 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4280 VDD.t1256 a_33497_n9032 a_34176_n6976 VDD.t1255 pfet_06v0 ad=0.3432p pd=2.44u as=0.2028p ps=1.3u w=0.78u l=0.5u
D119 a_21692_n6694.t29 VDD.t644 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X4281 VDD.t3422 a_39052_n12645 a_38964_n12548 VDD.t3421 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4282 a_13501_n22528.t11 a_11023_n22908.t38 a_11087_n23528.t15 VDD.t214 pfet_03v3 ad=1.82p pd=6.9u as=0.728p ps=3.32u w=2.8u l=0.28u
X4283 a_24964_n14116 a_24516_n14475 VDD.t3981 VDD.t3980 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X4284 a_46243_769 a_46573_841 a_46693_951 VSS.t2805 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X4285 a_32533_n12952 a_32413_n12996 a_31789_n12996 VSS.t932 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X4286 VDD.t2482 a_42972_n2804 a_42884_n2760 VDD.t2481 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4287 VDD.t684 a_13623_n6840.t41 a_11023_n6840.t18 VDD.t683 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4288 a_22444_332.t1 a_25836_n1236.t39 VDD.t3734 VDD.t3733 pfet_06v0 ad=0.2561p pd=1.505u as=0.30535p ps=1.605u w=0.985u l=0.5u
X4289 a_30180_n12168 a_21692_n6694.t30 a_29920_n12168 VDD.t645 pfet_06v0 ad=0.1736p pd=1.18u as=0.224p ps=1.36u w=0.56u l=0.5u
X4290 a_28940_n2406.t1 a_24631_n3588 VDD.t3221 VDD.t3220 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X4291 VSS.t3513 a_26060_n878.t3 a_25524_n708 VSS.t3512 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4292 a_29056_n14432 a_26944_n14116 a_28744_n14432 VDD.t3919 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X4293 a_13623_n22908.t6 a_21772_n452.t17 VSS.t1683 VSS.t1682 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4294 a_21792_n7464 a_21692_n7508.t3 VSS.t4342 VSS.t682 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X4295 VSS.t908 a_21772_n3588.t17 a_13623_n20230.t1 VSS.t907 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4296 VDD.t2179 a_39948_n6373 a_39860_n6276 VDD.t2178 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4297 VDD.t3350 a_25627_n452 a_25539_n407.t1 VDD.t3349 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X4298 VDD.t2377 a_24760_n11383 a_24672_n11339 VDD.t2376 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4299 VDD.t2947 a_39948_n3237 a_39860_n3140 VDD.t2946 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4300 a_28548_n5112 a_24815_n3588.t19 a_30884_n5112 VSS.t25 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X4301 VDD.t3399 a_41852_n7508 a_41764_n7464 VDD.t3398 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4302 a_13501_n19850.t11 a_13623_n20230.t41 a_11087_n20850.t21 VSS.t639 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4303 a_11087_n7460.t30 a_2167_3472.t81 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X4304 VDD.t3784 a_40956_n15348 a_40868_n15304 VDD.t3783 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D120 a_22220_690.t15 VDD.t783 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X4305 VDD.t1538 a_41852_n4372 a_41764_n4328 VDD.t1537 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D121 a_23072_n13432.t96 VDD.t533 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X4306 a_11087_n20850.t20 a_13623_n20230.t42 a_13501_n19850.t10 VSS.t640 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X4307 a_27337_1944.t0 a_26607_1966 VSS.t3755 VSS.t3754 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X4308 VDD.t647 a_21692_n6694.t31 a_29532_n4372.t1 VDD.t646 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4309 VDD.t3972 a_38716_n16916 a_38628_n16872 VDD.t3971 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4310 a_11023_n9518.t12 a_13623_n9518.t33 VDD.t268 VDD.t267 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4311 a_22588_n18917 a_22500_n18820 VSS.t1288 VSS.t1287 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4312 VDD.t4000 a_38716_n13780 a_38628_n13736 VDD.t3999 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4313 VDD.t566 a_13623_n4162.t42 a_11023_n4162.t12 VDD.t565 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4314 VSS.t3608 a_32543_n9032 a_33019_n8457 VSS.t3607 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X4315 VDD.t3831 a_36588_n18917 a_36500_n18820 VDD.t3830 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4316 VDD.t2586 a_24828_n20052 a_24740_n20008 VDD.t2585 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4317 a_11087_n15494.t33 a_2167_3472.t10 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X4318 a_13501_n22528.t1 a_13623_n22908.t34 a_11087_n23528.t1 VSS.t230 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4319 VDD.t2816 a_31772_n16916 a_31684_n16872 VDD.t2815 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4320 a_36924_n20485 a_36836_n20388 VSS.t1524 VSS.t1523 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4321 a_11087_n23528.t57 a_2167_3472.t45 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X4322 a_34796_n13780 a_34708_n13736 VSS.t2707 VSS.t2706 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4323 VDD.t359 a_21692_n5468.t30 a_21604_n708 VDD.t358 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X4324 a_27804_n14165 a_27496_n14116 VDD.t1978 VDD.t1977 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X4325 a_32543_n9032 a_31919_n9032 a_32395_n8456 VSS.t2220 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4326 a_35804_n20485 a_35716_n20388 VSS.t2054 VSS.t2053 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4327 VDD.t875 a_34348_n18917 a_34260_n18820 VDD.t874 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4328 OUT[0].t8 a_29408_1944.t23 VDD.t3910 VDD.t3909 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4329 VSS.t606 a_13623_n4162.t43 a_2167_3472.t9 VSS.t605 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4330 a_34544_n2272 a_32020_n2276 a_34232_n2272 VSS.t3106 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X4331 VSS.t3775 a_27337_1944.t3 a_22820_n2804 VSS.t3774 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X4332 VDD.t1023 a_24233_n8684 a_24128_n8544 VDD.t1022 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X4333 VDD.t1067 a_21916_n6694.t20 a_28852_n8292.t0 VDD.t1066 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X4334 a_38716_n20052 a_38628_n20008 VSS.t2277 VSS.t2276 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4335 VSS.t884 a_33776_n5896.t21 a_34708_n5896.t1 VSS.t883 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X4336 VSS.t2304 a_29900_760.t16 a_38996_n408 VSS.t2303 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4337 VDD.t2951 a_24233_n5548 a_24128_n5408 VDD.t2950 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X4338 VDD.t184 a_33496_n6659.t37 a_31628_n5940.t18 VDD.t183 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4339 a_11087_n23528.t58 a_2167_3472.t44 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X4340 EOC.t3 a_45648_1564.t19 VSS.t37 VSS.t36 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4341 a_28736_n4633.t15 a_30452_n5156.t13 a_30378_n5112 VSS.t1084 nfet_06v0 ad=0.4161p pd=1.905u as=0.1517p ps=1.19u w=0.82u l=0.6u
X4342 a_24233_n8684 a_23816_n8544 a_24609_n8544 VSS.t1767 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X4343 a_24569_n11820 a_24152_n11680 a_24945_n11680 VSS.t2998 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X4344 a_31772_n20052 a_31684_n20008 VSS.t2247 VSS.t2246 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4345 a_24233_n5548 a_23816_n5408 a_24609_n5408 VSS.t3117 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X4346 VDD.t1677 a_24752_n16132 a_23564_n8292 VDD.t1676 pfet_06v0 ad=0.35315p pd=1.96u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4347 a_26154_n4536 a_25530_n5112 a_25986_n4536 VDD.t3760 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X4348 VDD.t102 a_13623_n17552.t41 a_11023_n17552.t12 VDD.t101 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4349 a_30192_n15304.t3 a_27988_n20388 VDD.t2735 VDD.t2734 pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X4350 a_25559_n12548 a_26239_n12996 VDD.t3213 VDD.t3212 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4351 VDD.t456 a_21772_1116.t18 a_13623_n4162.t9 VDD.t455 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4352 a_13501_n6460.t4 a_13623_n6840.t42 a_11087_n7460.t7 VSS.t744 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4353 a_29532_n18484 a_29444_n18440 VSS.t2634 VSS.t2633 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4354 a_11023_n17552.t11 a_13623_n17552.t42 VDD.t104 VDD.t103 pfet_03v3 ad=0.728p pd=3.32u as=1.82p ps=6.9u w=2.8u l=0.28u
X4355 VDD.t3865 a_29900_n10600.t9 a_29532_n4372.t2 VDD.t3864 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4356 a_22352_n12097 a_21940_n11684 VSS.t2273 VSS.t2272 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4357 VDD.t2598 a_46108_n20052 a_46020_n20008 VDD.t2597 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4358 a_33280_n13248 a_31664_n13292 a_32152_n13692 VSS.t1811 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4359 a_42748_n4372 a_42660_n4328 VSS.t2735 VSS.t2734 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4360 a_28736_n4633.t10 a_30452_n5156.t14 VDD.t1049 VDD.t1048 pfet_06v0 ad=0.2197p pd=1.365u as=0.4056p ps=1.805u w=0.845u l=0.5u
X4361 a_10778_2852.t9 a_10712_4516.t51 VSS.t355 VSS.t354 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
D122 VSS.t4142 a_22140_n6694.t16 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X4362 VDD.t2362 a_43980_n11077 a_43892_n10980 VDD.t2361 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4363 VSS.t3054 a_34428_n452.t7 a_37396_1205 VSS.t3053 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4364 VSS.t4039 a_29211_n6724 a_29123_n6679 VSS.t4038 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X4365 VDD.t1758 a_13623_n12196.t43 a_11023_n12196.t18 VDD.t1757 pfet_03v3 ad=1.82p pd=6.9u as=0.728p ps=3.32u w=2.8u l=0.28u
X4366 VDD.t1558 a_46556_n18484 a_46468_n18440 VDD.t1557 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4367 VSS.t2376 a_30192_n15304.t21 a_24481_761.t5 VSS.t2375 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X4368 a_39164_n9076 a_39076_n9032 VSS.t1410 VSS.t1409 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4369 a_11023_n12196.t19 a_13623_n12196.t44 VDD.t1760 VDD.t1759 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4370 VSS.t4306 a_23564_n17700 a_21772_n17700.t0 VSS.t4305 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
D123 VSS.t695 a_21692_n6694.t32 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X4371 a_29127_n1400 a_28671_n1976 VDD.t3781 VDD.t3780 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X4372 a_33900_n17349 a_33812_n17252 VSS.t2695 VSS.t2694 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4373 a_13623_n9518.t0 a_21772_n17700.t23 VSS.t1057 VSS.t1056 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4374 a_24481_761.t7 a_30192_n15304.t22 VSS.t2378 VSS.t2377 nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X4375 VSS.t3816 a_23564_n14564.t9 a_21772_n14564.t0 VSS.t3815 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4376 VDD.t997 a_25237_n10599 a_25642_n9816 VDD.t996 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X4377 a_30136_n10600 a_29076_n8292.t10 VSS.t471 VSS.t470 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4378 VDD.t2490 a_41740_n11077 a_41652_n10980 VDD.t2489 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4379 VDD.t1706 a_25539_n407.t5 a_25759_1944 VDD.t1705 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X4380 a_25084_1564 a_24628_1252 VDD.t3629 VDD.t3628 pfet_06v0 ad=0.5368p pd=3.32u as=0.35315p ps=1.96u w=1.22u l=0.5u
X4381 a_28836_376 a_28132_376 VSS.t3771 VSS.t3770 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4382 VDD.t1866 a_44428_n9509 a_44340_n9412 VDD.t1865 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D124 a_25940_n17606.t23 VDD.t4122 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X4383 VSS.t2319 a_26755_n16132 a_26239_n12996 VSS.t2318 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4384 a_33900_n14213 a_33812_n14116 VSS.t4154 VSS.t4153 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4385 a_13623_n12196.t0 a_21772_n14564.t19 VSS.t1605 VSS.t1604 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4386 a_23816_n704 a_21604_n708 a_22876_n1148 VDD.t3357 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X4387 a_25879_n4328 a_25423_n4328 VDD.t1335 VDD.t1334 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X4388 VDD.t2494 a_40620_n11077 a_40532_n10980 VDD.t2493 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4389 VDD.t1316 a_13623_n14874.t42 a_11023_n14874.t17 VDD.t1315 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4390 VSS.t894 a_4001_4292.t11 a_10778_2852.t14 VSS.t336 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4391 a_25948_n20485 a_25860_n20388 VSS.t4082 VSS.t4081 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4392 a_11023_n14874.t18 a_13623_n14874.t43 VDD.t1318 VDD.t1317 pfet_03v3 ad=0.728p pd=3.32u as=1.82p ps=6.9u w=2.8u l=0.28u
X4393 VSS.t2572 a_44004_n1192 a_44640_1944.t0 VSS.t2571 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4394 VSS.t2768 a_11023_n4162.t38 VSS.t2768 VSS.t54 nfet_03v3 ad=0.728p pd=3.32u as=0 ps=0 w=2.8u l=0.28u
X4395 VDD.t824 a_34708_n5896.t28 a_33496_n8222.t3 VDD.t823 pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X4396 a_26692_1564 a_25524_1243 a_26488_1564 VDD.t1364 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X4397 VDD.t2302 a_39164_n12212 a_39076_n12168 VDD.t2301 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4398 a_28736_n4633.t0 a_24815_n3588.t20 VDD.t38 VDD.t37 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X4399 VDD.t3500 a_35064_n11383 a_28300_n15348 VDD.t3499 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4400 a_26563_n12212 a_21996_n12996.t12 a_27524_n15304 VDD.t3490 pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4401 VSS.t910 a_21772_n3588.t18 a_13623_n20230.t0 VSS.t909 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4402 VDD.t4256 a_25500_n20485 a_25412_n20388 VDD.t4255 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4403 a_23619_n9860 a_23949_n9860 a_24069_n9262 VDD.t1930 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X4404 a_24935_n3544 a_24815_n3588.t21 a_24751_n3544 VSS.t26 nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X4405 a_27337_n3140 a_26607_n3544 VDD.t4235 VDD.t4234 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X4406 a_23619_n6724 a_23949_n6724 a_24069_n6126 VDD.t920 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X4407 a_44004_n1192 a_43556_n661 VDD.t1331 VDD.t1330 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X4408 a_38604_n12645 a_38516_n12548 VSS.t2158 VSS.t2157 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4409 a_42476_1515 a_42168_1564 VSS.t1810 VSS.t1809 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X4410 a_11023_n22908.t11 a_13623_n22908.t35 VDD.t233 VDD.t232 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4411 VDD.t2945 a_43196_n16916 a_43108_n16872 VDD.t2944 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4412 a_32984_n2672 a_32432_n2689 a_32780_n2672 VDD.t3388 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X4413 a_45324_n7941 a_45236_n7844 VSS.t1470 VSS.t1469 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4414 a_23816_n704 a_22016_n1121 a_22876_n1148 VSS.t3438 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X4415 VDD.t235 a_13623_n22908.t36 a_11023_n22908.t10 VDD.t234 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4416 VDD.t3537 a_43196_n13780 a_43108_n13736 VDD.t3536 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4417 VDD.t346 a_10712_4516.t52 a_10778_2852.t1 VDD.t345 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4418 a_26839_n2990 a_26383_n2968 a_26607_n3544 VDD.t1613 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X4419 a_29612_n8292 a_28736_n4633.t23 VDD.t1037 VDD.t1036 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X4420 a_47228_n20485 a_47140_n20388 VSS.t1065 VSS.t1064 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4421 VSS.t2693 a_26328_n6654.t22 a_21692_n13308.t0 VSS.t2692 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X4422 VDD.t849 a_25020_n8200.t7 a_29532_n10311 VDD.t848 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4423 a_43196_n9076 a_43108_n9032 VSS.t3186 VSS.t3185 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D125 VSS.t825 a_24481_761.t91 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X4424 VSS.t921 a_40652_n1572 a_45648_1564.t0 VSS.t920 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4425 VDD.t3133 a_45212_n5940 a_45124_n5896 VDD.t3132 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4426 VSS.t3805 a_25836_n1236.t40 a_24631_n3588 VSS.t3804 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X4427 VDD.t2278 a_38828_n11077 a_38740_n10980 VDD.t2277 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4428 a_45648_1564.t5 a_40652_n1572 VDD.t869 VDD.t868 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4429 VDD.t4289 a_45212_n2804 a_45124_n2760 VDD.t4288 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4430 a_34552_n3140 a_33588_n3461 a_34348_n3140 VSS.t3419 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4431 a_27167_n10808 a_26543_n11384 a_26999_n10808 VDD.t1947 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X4432 a_31909_n12398 a_31789_n12996 VDD.t4298 VDD.t4297 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X4433 VDD.t202 a_38256_1564.t22 OUT[3].t9 VDD.t201 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4434 a_43196_n20052 a_43108_n20008 VSS.t3896 VSS.t3895 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4435 VDD.t3107 a_23703_n5156.t9 a_25559_n12548 VDD.t3106 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4436 a_11087_n23528.t59 a_2167_3472.t43 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X4437 a_27348_n2672 a_25547_n2445 a_26499_n2732 VDD.t3891 pfet_06v0 ad=0.1313p pd=1.025u as=0.19315p ps=1.27u w=0.505u l=0.5u
X4438 VDD.t186 a_33496_n6659.t38 a_31628_n5940.t17 VDD.t185 pfet_06v0 ad=0.428p pd=2.02u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4439 a_22364_n13648 a_22264_n13692 VSS.t1607 VSS.t1606 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4440 a_28009_n1192.t1 a_27279_n1170 VDD.t2118 VDD.t2117 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X4441 a_35848_n3868 a_25237_n4327 VSS.t1206 VSS.t1205 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X4442 a_22892_n5156.t0 a_30555_n2729 a_32132_n4708 VDD.t2978 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X4443 a_13501_n19850.t0 a_11023_n20230.t38 a_11087_n20850.t18 VDD.t1905 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4444 a_25627_n452 a_25975_n184 VDD.t1353 VDD.t1352 pfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X4445 a_45212_n9076 a_45124_n9032 VSS.t3663 VSS.t3662 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4446 a_23932_n18917 a_23844_n18820 VSS.t3646 VSS.t1942 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4447 VDD.t1200 a_38403_n5503 a_36773_n5468 VDD.t1199 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4448 a_43728_1248 a_41204_1243 a_43416_1248 VSS.t1867 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X4449 a_38295_332 a_38951_420 a_38847_464 VDD.t3216 pfet_06v0 ad=0.25375p pd=1.51u as=0.1313p ps=1.025u w=0.505u l=0.5u
X4450 VSS.t2501 a_23999_n2320.t7 a_25647_n1976 VSS.t2500 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X4451 a_32308_n1976 a_29076_n8292.t11 a_32308_n1572 VDD.t442 pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4452 a_33538_n12168 a_32854_n12168 VDD.t2858 VDD.t2857 pfet_06v0 ad=61.199993f pd=0.7u as=0.1656p ps=1.28u w=0.36u l=0.5u
X4453 VDD.t1438 a_37932_n18917 a_37844_n18820 VDD.t1437 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4454 VDD.t1389 a_39724_n17349 a_39636_n17252 VDD.t1388 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4455 a_29161_n14476 a_28744_n14432 a_29537_n14432 VSS.t2627 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X4456 VDD.t1450 a_38403_n2367 a_37452_n3888 VDD.t1449 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4457 a_11023_n9518.t0 a_13623_n9518.t34 VSS.t267 VSS.t266 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4458 a_47564_n17349 a_47476_n17252 VSS.t3887 VSS.t3886 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4459 VDD.t1713 a_37368_n320 a_37785_n364 VDD.t1712 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X4460 a_27511_n12146 a_27055_n12168 a_27279_n12146 VDD.t2853 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X4461 VDD.t940 a_39724_n14213 a_39636_n14116 VDD.t939 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4462 a_21772_n452.t1 a_23564_n452.t8 VDD.t3664 VDD.t3663 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4463 a_24128_n3840 a_22016_n4257 a_23816_n3840 VDD.t3264 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X4464 a_27042_n4536 a_26358_n4618 VDD.t1400 VDD.t1399 pfet_06v0 ad=61.199993f pd=0.7u as=0.1656p ps=1.28u w=0.36u l=0.5u
X4465 a_11023_n20230.t11 a_13623_n20230.t43 VDD.t594 VDD.t593 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4466 a_47564_n14213 a_47476_n14116 VSS.t3555 VSS.t3554 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4467 a_24693_n9240 a_24573_n9860 a_23949_n9860 VDD.t996 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X4468 a_22904_n12080 a_22352_n12097 a_22700_n12080 VDD.t0 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
D126 VSS.t14 a_22444_332.t33 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X4469 VSS.t550 a_23072_n13432.t97 a_23024_n8544 VSS.t549 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4470 VDD.t596 a_13623_n20230.t44 a_11023_n20230.t10 VDD.t595 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4471 a_45324_n17349 a_45236_n17252 VSS.t3190 VSS.t3189 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4472 VDD.t924 a_31660_n17349 a_31572_n17252 VDD.t923 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4473 a_27055_n1192 a_26431_n1192 a_26887_n1192 VDD.t3189 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X4474 VSS.t3677 a_23004_n2332 a_22940_n2276 VSS.t3676 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X4475 a_45324_n14213 a_45236_n14116 VSS.t3192 VSS.t3191 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4476 a_33216_1944.t4 a_25084_1564 VDD.t1123 VDD.t1122 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4477 VSS.t552 a_23072_n13432.t98 a_23024_n5408 VSS.t551 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4478 a_36709_n5412 a_28736_n4633.t24 VSS.t1074 VSS.t1073 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4479 a_13623_n4162.t8 a_21772_1116.t19 VDD.t460 VDD.t459 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4480 a_11023_n4162.t11 a_13623_n4162.t44 VDD.t568 VDD.t567 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4481 a_31076_376 a_30372_376 VDD.t3932 VDD.t3931 pfet_06v0 ad=0.3477p pd=1.79u as=0.4392p ps=1.94u w=1.22u l=0.5u
X4482 VDD.t2584 a_44876_n9509 a_44788_n9412 VDD.t2583 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4483 VSS.t71 a_11023_n14874.t37 a_11087_n15494.t21 VSS.t70 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4484 VDD.t361 a_21692_n5468.t31 a_29444_n708 VDD.t360 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X4485 VDD.t1232 a_41852_n10644 a_41764_n10600 VDD.t1231 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4486 a_27524_n15304 a_27404_n14990 VDD.t3274 VDD.t3273 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
D127 VSS.t1314 a_21804_n2273.t13 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X4487 VDD.t2965 a_33608_n4284 a_33416_n4240 VDD.t2964 pfet_06v0 ad=0.2222p pd=1.89u as=0.2424p ps=1.465u w=0.505u l=0.5u
X4488 VDD.t3312 a_37372_n9076 a_37284_n9032 VDD.t3311 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4489 a_11087_n15494.t20 a_11023_n14874.t38 VSS.t73 VSS.t72 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X4490 VDD.t987 a_39164_n20485 a_39076_n20388 VDD.t986 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4491 VDD.t1244 a_36812_n7941 a_36724_n7844 VDD.t1243 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4492 a_11087_n10138.t16 a_11023_n9518.t36 a_13501_n9138.t8 VDD.t549 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4493 a_33686_n11592 a_32854_n12168 a_33518_n11592 VSS.t2921 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4494 a_30864_n704 a_30716_n1148 a_30696_n704 VSS.t1999 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4495 a_22940_n2276 a_22820_n2804 a_22672_n2214.t2 VSS.t3948 nfet_06v0 ad=0.1312p pd=1.14u as=0.2569p ps=1.56u w=0.82u l=0.6u
X4496 a_28644_n9815 a_26388_n17606.t11 a_28624_n9394 VSS.t366 nfet_06v0 ad=0.2119p pd=1.335u as=0.4137p ps=1.9u w=0.815u l=0.6u
X4497 VDD.t2227 a_29900_760.t17 a_41684_n1976 VDD.t2226 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4498 a_39477_n2184 a_39357_n2228 a_38733_n2295 VSS.t2838 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X4499 VSS.t4088 a_31961_n11340 a_31856_n11296 VSS.t4087 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X4500 a_30584_1248 a_29744_1564 a_30296_1564 VSS.t1157 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4501 VDD.t1574 a_43416_1248 a_43833_1204 VDD.t1573 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X4502 a_41852_n16916 a_41764_n16872 VSS.t2132 VSS.t2131 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4503 a_33292_n2716 a_32984_n2672 VDD.t1972 VDD.t1971 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X4504 VDD.t2383 a_24264_n6976 a_24681_n7116 VDD.t2382 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X4505 VSS.t3942 a_24573_n9860 a_24693_n9816 VSS.t3941 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4506 VDD.t1472 a_47900_n18484 a_47812_n18440 VDD.t1471 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4507 a_23823_n5111 a_23703_n5156.t10 a_23228_n6679 VSS.t3183 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X4508 a_35456_n4628.t3 a_34708_n5896.t29 VDD.t826 VDD.t825 pfet_06v0 ad=0.2952p pd=1.54u as=0.3608p ps=2.52u w=0.82u l=0.5u
X4509 VSS.t2362 a_21812_n6643 a_25412_n8501 VSS.t2361 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4510 a_43084_n12645 a_42996_n12548 VSS.t1482 VSS.t1481 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4511 a_11087_n7460.t8 a_13623_n6840.t43 a_13501_n6460.t1 VSS.t745 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4512 VSS.t1076 a_28736_n4633.t25 a_29476_n6980 VSS.t1075 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4513 VSS.t124 a_11023_n12196.t37 a_11087_n12816.t1 VSS.t70 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4514 VDD.t3521 a_29868_n17349 a_29780_n17252 VDD.t3520 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4515 a_45772_n7941 a_45684_n7844 VSS.t3536 VSS.t3535 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4516 VDD.t1442 a_26956_n18917 a_26868_n18820 VDD.t1441 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4517 a_11087_n18172.t20 a_11023_n17552.t38 VSS.t419 VSS.t56 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4518 a_11087_n12816.t0 a_11023_n12196.t38 VSS.t125 VSS.t72 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X4519 VSS.t2011 a_37859_377 a_39748_2475 VSS.t2010 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4520 a_27988_n4328 a_27540_n3797 VSS.t2267 VSS.t2266 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X4521 a_13501_n9138.t10 a_13623_n9518.t35 a_11087_n10138.t27 VSS.t268 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4522 a_36588_n17349 a_36500_n17252 VSS.t2605 VSS.t2604 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4523 a_25972_n6276 a_25524_n6635 VDD.t3300 VDD.t3299 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X4524 a_30320_n6636 a_31548_n10172.t24 VSS.t290 VSS.t289 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4525 a_36588_n14213 a_36500_n14116 VSS.t4213 VSS.t4212 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4526 VDD.t1509 a_33077_n1191 a_35940_n1931 VDD.t1508 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X4527 VDD.t3251 a_45660_n5940 a_45572_n5896 VDD.t3250 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4528 a_34348_n17349 a_34260_n17252 VSS.t2608 VSS.t2607 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4529 a_30612_n1104 a_29444_n708 a_30408_n1104 VDD.t2742 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X4530 VDD.t2026 a_45660_n2804 a_45572_n2760 VDD.t2025 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4531 VDD.t4097 a_42188_n11077 a_42100_n10980 VDD.t4096 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4532 VDD.t3124 a_28752_n15348 a_28212_n15303 VDD.t3123 pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X4533 a_34348_n14213 a_34260_n14116 VSS.t3890 VSS.t2256 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4534 VSS.t2078 CLK.t14 a_33496_n6659.t7 VSS.t2077 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4535 VSS.t2809 a_27988_n20388 a_30192_n15304.t0 VSS.t2808 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4536 a_46556_n12212 a_46468_n12168 VSS.t3620 VSS.t3619 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4537 a_11087_n10138.t31 a_2167_3472.t82 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X4538 a_32108_n17349 a_32020_n17252 VSS.t3892 VSS.t3891 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4539 a_30472_n9815 a_28617_n8548 VSS.t2650 VSS.t2649 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X4540 a_34652_n11391 a_34089_n10252 VDD.t1518 VDD.t1517 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X4541 VSS.t1691 a_30732_332.t7 a_35940_2475 VSS.t1690 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4542 VSS.t1329 a_27672_n3543 a_21692_n7508.t0 VSS.t1328 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X4543 VDD.t785 a_22220_690.t16 a_37585_n3140 VDD.t784 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X4544 VDD.t2899 a_44540_n7508 a_44452_n7464 VDD.t2898 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4545 VDD.t2193 a_38716_n20052 a_38628_n20008 VDD.t2192 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4546 a_11087_n20850.t19 a_11023_n20230.t39 VSS.t1979 VSS.t58 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4547 VDD.t3042 a_45660_n16916 a_45572_n16872 VDD.t3041 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4548 EOC.t2 a_45648_1564.t20 VSS.t39 VSS.t38 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4549 VSS.t848 a_25612_n878.t7 a_21916_n1975 VSS.t847 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X4550 VDD.t2276 a_44540_n16916 a_44452_n16872 VDD.t2275 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4551 VDD.t3532 a_44540_n4372 a_44452_n4328 VDD.t3531 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4552 a_45660_n9076 a_45572_n9032 VSS.t1339 VSS.t1338 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4553 VDD.t3666 a_45660_n13780 a_45572_n13736 VDD.t3665 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4554 VDD.t3215 a_41336_n407 a_24236_2258.t1 VDD.t3214 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4555 a_34455_n1422 a_33999_n1400 a_34223_n1976 VDD.t3443 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X4556 a_22700_n12080 a_22600_n12124 VDD.t1549 VDD.t1548 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X4557 VDD.t2167 a_31772_n20052 a_31684_n20008 VDD.t2166 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4558 VDD.t2126 a_44540_n13780 a_44452_n13736 VDD.t2125 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4559 VDD.t3512 a_32860_n2020 a_32736_n1572 VDD.t3511 pfet_06v0 ad=0.6588p pd=3.52u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4560 a_21892_n12952 a_22220_n12996 a_21872_n12530 VSS.t4281 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4561 VDD.t1901 a_47116_n18917 a_47028_n18820 VDD.t1900 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4562 VSS.t357 a_10712_4516.t53 a_10778_2852.t2 VSS.t356 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4563 a_30244_860 a_28492_332 VSS.t1412 VSS.t1411 nfet_06v0 ad=0.1968p pd=1.3u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4564 a_28841_n3844 a_28144_n4708 a_27932_n3543 VSS.t3830 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X4565 VDD.t3179 a_42300_n16916 a_42212_n16872 VDD.t3178 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4566 a_24576_n6976 a_22464_n7393 a_24264_n6976 VDD.t4044 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X4567 VDD.t1137 a_41292_n18917 a_41204_n18820 VDD.t1136 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4568 VDD.t1833 a_43084_n17349 a_42996_n17252 VDD.t1832 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4569 a_26702_n13736 a_26266_n13736 a_26470_n13736 VDD.t4257 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X4570 a_47317_376 a_47197_908 a_46573_841 VDD.t2649 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X4571 a_33608_n4284 a_33015_n4284 a_34344_n3840 VSS.t2878 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4572 a_30876_n16916 a_30788_n16872 VSS.t4274 VSS.t4273 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4573 VDD.t3452 a_42300_n13780 a_42212_n13736 VDD.t3451 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4574 a_26736_n364 a_21692_n5468.t32 VDD.t363 VDD.t362 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
D128 VSS.t15 a_22444_332.t34 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X4575 a_26328_n6654.t0 a_28156_n6412.t29 VSS.t712 VSS.t711 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4576 a_22700_n12080 a_22600_n12124 VSS.t1626 VSS.t1625 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4577 VDD.t1540 a_40172_n18917 a_40084_n18820 VDD.t1539 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4578 VDD.t1909 a_25160_n14816 a_25577_n14956 VDD.t1908 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X4579 VDD.t4012 a_43084_n14213 a_42996_n14116 VDD.t4011 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4580 VSS.t3362 a_26172_n14564.t3 a_25636_n14520 VSS.t3361 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4581 a_11087_n15494.t10 a_11023_n14874.t39 a_13501_n14494.t10 VDD.t82 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4582 VDD.t2443 a_47116_n101 a_47028_n4 VDD.t2442 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4583 a_45660_n20052 a_45572_n20008 VSS.t3971 VSS.t3970 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4584 VDD.t1946 a_35804_n18484 a_35716_n18440 VDD.t1945 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4585 a_11023_n9518.t11 a_13623_n9518.t36 VDD.t270 VDD.t269 pfet_03v3 ad=0.728p pd=3.32u as=1.82p ps=6.9u w=2.8u l=0.28u
X4586 a_44540_n20052 a_44452_n20008 VSS.t3975 VSS.t3974 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4587 a_30204_n1104 a_30104_n1148 VDD.t4029 VDD.t4028 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X4588 VDD.t1484 a_29295_n1400 a_29751_n1422 VDD.t1483 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X4589 a_22164_n2760 a_21716_n2229 VDD.t3994 VDD.t3993 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X4590 a_40172_n9509 a_40084_n9412 VSS.t2616 VSS.t2615 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4591 a_31872_n10529 a_31460_n10116 VDD.t1277 VDD.t1276 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X4592 a_10778_2852.t14 a_4001_4292.t12 VSS.t895 VSS.t338 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X4593 a_41740_n6373 a_41652_n6276 VSS.t2619 VSS.t2618 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4594 a_42300_n20052 a_42212_n20008 VSS.t4341 VSS.t4340 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4595 a_26060_n18917 a_25972_n18820 VSS.t974 VSS.t973 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4596 a_11087_n18172.t10 a_11023_n17552.t39 a_13501_n17172.t10 VDD.t409 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4597 a_33494_n9860 a_28519_n10160.t9 VDD.t791 VDD.t790 pfet_06v0 ad=0.5368p pd=3.32u as=0.4941p ps=2.03u w=1.22u l=0.5u
X4598 a_33467_1116 a_33815_1384 VDD.t1001 VDD.t1000 pfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X4599 a_44428_n4805 a_44340_n4708 VSS.t1567 VSS.t1566 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4600 a_22568_n13648 a_21604_n13252 a_22364_n13648 VSS.t2216 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4601 VDD.t535 a_23072_n13432.t99 a_32412_n13648 VDD.t534 pfet_06v0 ad=0.45p pd=2.02u as=0.3432p ps=2.44u w=0.78u l=0.5u
X4602 VSS.t138 a_31628_n5940.t43 a_33776_n5896.t1 VSS.t137 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4603 VDD.t433 a_33216_1944.t22 OUT[1].t9 VDD.t432 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4604 a_43868_n2804 a_43780_n2760 VSS.t2401 VSS.t2400 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4605 VDD.t1355 a_46668_n6373 a_46580_n6276 VDD.t1354 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4606 a_22568_n8944 a_21604_n8548 a_22364_n8944 VSS.t4030 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4607 a_11087_n12816.t10 a_11023_n12196.t39 a_13501_n11816.t0 VDD.t136 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4608 VDD.t3004 a_42748_n15348 a_42660_n15304 VDD.t3003 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4609 VDD.t3837 a_46668_n3237 a_46580_n3140 VDD.t3836 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4610 a_28433_n3844 a_27337_n3140 VSS.t3105 VSS.t3104 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X4611 a_22568_n5808 a_21604_n5412 a_22364_n5808 VSS.t3578 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4612 a_28212_n15303 a_21692_n6694.t33 a_27404_n14990 VDD.t648 pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4613 a_11087_n15494.t9 a_13623_n14874.t44 a_13501_n14494.t9 VSS.t1373 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4614 a_26719_n7464 a_26095_n7464 a_26571_n6888 VSS.t1159 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4615 VDD.t2477 a_40508_n15348 a_40420_n15304 VDD.t2476 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4616 a_39352_464 a_39056_820 a_38295_332 VDD.t945 pfet_06v0 ad=0.2424p pd=1.465u as=0.25375p ps=1.51u w=0.505u l=0.5u
X4617 VSS.t1510 a_38403_n2367 a_37452_n3888 VSS.t1509 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4618 VDD.t2633 a_21692_n13308.t33 a_21604_n8548 VDD.t2632 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X4619 a_35064_n11383 a_34350_n10980 VDD.t1466 VDD.t1465 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X4620 VDD.t3035 a_33564_n16916 a_33476_n16872 VDD.t3034 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4621 VSS.t278 a_44640_1944.t22 OUT[5].t1 VSS.t277 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4622 VDD.t365 a_21692_n5468.t33 a_21604_n5412 VDD.t364 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X4623 a_13501_n17172.t1 a_13623_n17552.t43 a_11087_n18172.t1 VSS.t102 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4624 a_43221_398 a_43101_841 VDD.t1849 VDD.t1848 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X4625 a_38716_n20485 a_38628_n20388 VSS.t4175 VSS.t4174 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4626 a_34796_n15348 a_34708_n15304 VSS.t2774 VSS.t1475 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4627 a_36588_n13780 a_36500_n13736 VSS.t2411 VSS.t2410 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4628 a_11087_n18172.t0 a_13623_n17552.t44 a_13501_n17172.t0 VSS.t103 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X4629 VDD.t1915 a_47116_n9509 a_47028_n9412 VDD.t1914 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4630 VDD.t3101 a_31324_n16916 a_31236_n16872 VDD.t3100 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4631 VDD.t3763 a_35692_n15348 a_35604_n15304 VDD.t2366 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4632 a_30652_n20485 a_30564_n20388 VSS.t1583 VSS.t1582 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4633 a_27224_n62 a_26736_n364 a_27484_n4 VDD.t1467 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X4634 VSS.t2126 a_29532_n4372.t8 a_30866_n3844 VSS.t2125 nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
X4635 a_27190_n5112 a_26358_n4618 a_27042_n4536 VDD.t1398 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X4636 VDD.t300 a_33496_n8222.t21 a_31548_n10172.t8 VDD.t299 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X4637 a_30871_n11728 a_33910_n12146 VDD.t3535 VDD.t3534 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X4638 a_23136_447 a_22724_860.t7 VDD.t863 VDD.t862 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
D129 a_25940_n17606.t24 VDD.t529 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X4639 a_33564_n20052 a_33476_n20008 VSS.t1758 VSS.t1757 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4640 VDD.t1585 a_24828_n18484 a_24740_n18440 VDD.t1584 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4641 a_11087_n12816.t29 a_13623_n12196.t45 a_13501_n11816.t19 VSS.t1849 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4642 a_33488_n12996 a_28927_n10160 VSS.t2393 VSS.t1813 nfet_06v0 ad=0.1584p pd=1.6u as=0.2344p ps=1.56u w=0.36u l=0.6u
X4643 VDD.t3145 a_33452_n15348 a_33364_n15304 VDD.t3144 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D130 a_22444_332.t35 VDD.t19 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X4644 a_10778_2852.t13 a_4001_4292.t13 VSS.t896 VSS.t340 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4645 a_27032_51 a_26631_7 a_25975_n184 VSS.t1487 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X4646 VSS.t1685 a_21772_n452.t18 a_13623_n22908.t7 VSS.t1684 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4647 a_31324_n20052 a_31236_n20008 VSS.t1237 VSS.t1236 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4648 a_28455_n10116 a_28335_n10644 VSS.t1131 VSS.t1130 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X4649 VSS.t3321 a_23619_n12996 a_22264_n13692 VSS.t3320 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4650 VDD.t3814 a_43196_n20052 a_43108_n20008 VDD.t3813 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4651 a_13501_n22528.t10 a_11023_n22908.t39 a_11087_n23528.t14 VDD.t215 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4652 VDD.t2000 CLK.t15 a_33496_n6659.t5 VDD.t1999 pfet_06v0 ad=0.3608p pd=2.52u as=0.2542p ps=1.44u w=0.82u l=0.5u
X4653 a_23708_n15216 a_23608_n15260 VDD.t3310 VDD.t3309 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X4654 a_45648_1564.t4 a_40652_n1572 VDD.t867 VDD.t866 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4655 a_13501_n9138.t9 a_11023_n9518.t37 a_11087_n10138.t17 VDD.t550 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4656 VDD.t314 a_21772_n11428.t22 a_13623_n14874.t9 VDD.t313 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4657 a_24380_n18484 a_24292_n18440 VSS.t1693 VSS.t1692 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4658 VSS.t2769 a_11023_n4162.t39 a_2167_3472.t40 VDD.t2700 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4659 a_48012_n7941 a_47924_n7844 VSS.t2593 VSS.t2592 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4660 a_13623_n14874.t8 a_21772_n11428.t23 VDD.t316 VDD.t315 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4661 a_28300_n20485 a_28212_n20388 VSS.t4084 VSS.t4083 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4662 a_37932_n17349 a_37844_n17252 VSS.t2658 VSS.t2657 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D131 VSS.t826 a_24481_761.t92 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X4663 VDD.t2668 a_45772_n11077 a_45684_n10980 VDD.t2667 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4664 a_26299_n16388 a_25831_n12996 a_21772_n12996 VSS.t2611 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4665 a_22276_n1572.t0 a_21828_n1931 VSS.t3909 VSS.t3908 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X4666 a_23816_n8544 a_21604_n8548 a_22876_n8988 VDD.t3951 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X4667 a_22140_n18484 a_22052_n18440 VSS.t1695 VSS.t1694 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4668 a_23360_n15233 a_22948_n14820 VSS.t2107 VSS.t2106 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4669 a_37932_n14213 a_37844_n14116 VSS.t2697 VSS.t2696 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4670 a_10712_4516.t11 a_10778_2852.t31 VSS.t389 VSS.t388 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4671 a_22116_860 a_21996_332.t3 VSS.t465 VSS.t464 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4672 a_27597_n8292 a_24716_n5156.t7 VSS.t1380 VSS.t1379 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4673 a_30204_n1104 a_30104_n1148 VSS.t4105 VSS.t4104 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4674 a_23816_n5408 a_21604_n5412 a_22876_n5852 VDD.t3493 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X4675 VDD.t2670 a_43532_n11077 a_43444_n10980 VDD.t2669 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4676 a_22140_n15348 a_22052_n15304 VSS.t1273 VSS.t1272 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4677 a_11087_n23528.t60 a_2167_3472.t42 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X4678 VDD.t3120 a_46108_n18484 a_46020_n18440 VDD.t3119 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4679 a_26118_n13160 a_25642_n13736 VSS.t1230 VSS.t1229 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4680 a_32337_1248 a_24481_761.t93 VSS.t828 VSS.t827 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X4681 VSS.t41 a_45648_1564.t21 EOC.t1 VSS.t40 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
D132 VSS.t4197 a_25940_n17606.t25 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X4682 a_40172_n5940 a_40084_n5896 VSS.t4027 VSS.t4026 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4683 a_47900_n12212 a_47812_n12168 VSS.t3679 VSS.t3678 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4684 VDD.t2885 a_22588_n16916 a_22500_n16872 VDD.t2884 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4685 a_13501_n6460.t6 a_11023_n6840.t38 a_11087_n7460.t20 VDD.t116 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4686 VDD.t3048 a_31544_n11296 a_31961_n11340 VDD.t3047 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X4687 a_11087_n23528.t0 a_13623_n22908.t37 a_13501_n22528.t0 VSS.t231 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
D133 a_26388_n17606.t12 VDD.t351 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X4688 VDD.t2058 a_26635_n12996 a_26547_n12951 VDD.t2057 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X4689 a_31961_1204 a_31544_1248 a_32337_1248 VSS.t1299 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X4690 VDD.t616 a_29920_n3900.t21 a_28940_n2406.t1 VDD.t615 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X4691 a_21812_n6643 a_22140_n6694.t17 a_22016_n6276 VDD.t4065 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4692 a_29900_760.t0 a_33252_n1192 VSS.t1319 VSS.t1318 nfet_06v0 ad=0.2132p pd=1.34u as=0.2911p ps=1.53u w=0.82u l=0.6u
X4693 a_44876_n4805 a_44788_n4708 VSS.t2192 VSS.t2191 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4694 VSS.t3347 a_31405_n452 a_31525_n408 VSS.t3346 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4695 VSS.t3319 a_24731_n3124.t5 a_40299_n2276 VSS.t3318 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X4696 a_29076_n8292.t3 a_25019_n3588.t9 VDD.t3395 VDD.t3394 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4697 a_33048_n7420 a_32455_n7420 a_33784_n6976 VSS.t4319 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4698 a_27404_n14990 a_28300_n15348 a_28212_n15303 VDD.t2257 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X4699 a_22052_1944 a_21604_2475 VDD.t2294 VDD.t2293 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X4700 VDD.t650 a_21692_n6694.t34 a_34986_n9032 VDD.t649 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X4701 OUT[2].t8 a_37024_1944.t23 VDD.t2602 VDD.t2601 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4702 a_32262_n452 a_22444_332.t36 VDD.t21 VDD.t20 pfet_06v0 ad=0.5368p pd=3.32u as=0.4941p ps=2.03u w=1.22u l=0.5u
X4703 a_22588_n20052 a_22500_n20008 VSS.t1455 VSS.t1287 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4704 a_36217_n3500 a_35800_n3456 a_36593_n3456 VSS.t1628 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X4705 a_21772_1116.t3 a_23564_1116.t8 VDD.t3411 VDD.t2340 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4706 a_24152_n11680 a_21940_n11684 a_23212_n12124 VDD.t2188 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X4707 VSS.t3699 a_31459_n14564 a_30159_n13296 VSS.t3698 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4708 OUT[4].t0 a_41392_1944.t23 VSS.t1442 VSS.t1441 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4709 a_26527_51 a_25627_n452 VDD.t3348 VDD.t3347 pfet_06v0 ad=0.1313p pd=1.025u as=0.29465p ps=1.74u w=0.505u l=0.5u
X4710 a_28583_n3140 a_28736_1944 a_27452_n2716 VDD.t1230 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X4711 a_21892_n9816 a_21772_n9860 VSS.t2814 VSS.t2813 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4712 a_34572_n12645 a_34484_n12548 VSS.t2386 VSS.t2385 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4713 a_33776_n5896.t0 a_31628_n5940.t44 VSS.t140 VSS.t139 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X4714 a_11023_n6840.t19 a_13623_n6840.t44 VDD.t686 VDD.t685 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4715 VSS.t3541 a_26266_n9240 a_26742_n9816 VSS.t3540 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X4716 a_11087_n20850.t41 a_2167_3472.t29 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X4717 VDD.t106 a_13623_n17552.t45 a_11023_n17552.t10 VDD.t105 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4718 a_26175_n12951 a_23703_n5156.t11 a_25132_n16432 VSS.t3184 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X4719 a_29444_n4328.t0 a_27259_804.t16 a_30040_n3844 VSS.t857 nfet_06v0 ad=0.2132p pd=1.34u as=0.1722p ps=1.24u w=0.82u l=0.6u
X4720 VDD.t383 a_10778_2852.t32 a_10712_4516.t21 VDD.t382 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4721 a_10712_4516.t10 a_10778_2852.t33 VSS.t391 VSS.t390 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4722 a_34872_1619 a_34471_1575 a_33815_1384 VSS.t4036 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X4723 VDD.t3800 a_47564_n9509 a_47476_n9412 VDD.t3799 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4724 a_42076_n20485 a_41988_n20388 VSS.t4054 VSS.t4053 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4725 a_32581_n9860 a_29444_n4328.t9 a_33572_n10980 VDD.t1497 pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4726 VDD.t3069 a_44316_n1669 a_44228_n1572 VDD.t3068 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4727 a_47900_n4372 a_47812_n4328 VSS.t2226 VSS.t2225 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4728 a_29532_n4372.t0 a_21692_n6694.t35 VDD.t652 VDD.t651 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X4729 VDD.t1404 a_26547_n12951 a_26543_n11384 VDD.t1403 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
D134 a_23072_n13432.t100 VDD.t536 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X4730 VSS.t113 a_11023_n6840.t39 a_11087_n7460.t10 VSS.t64 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X4731 a_31544_n11296 a_29332_n11301 a_30604_n11029 VDD.t3473 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X4732 a_29076_n8292.t1 a_25836_n1236.t41 VDD.t3736 VDD.t3735 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X4733 VDD.t2875 a_39500_n7941 a_39412_n7844 VDD.t2874 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4734 a_26531_n8639 a_26861_n8567 a_26981_n8457 VSS.t3001 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X4735 a_41964_1564 a_41864_1394 VDD.t3880 VDD.t3879 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X4736 VDD.t40 a_24815_n3588.t22 a_34736_n3840 VDD.t39 pfet_06v0 ad=0.3432p pd=2.44u as=0.2028p ps=1.3u w=0.78u l=0.5u
X4737 VDD.t272 a_13623_n9518.t37 a_11023_n9518.t10 VDD.t271 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4738 a_38380_n15781 a_38292_n15684 VSS.t3562 VSS.t3561 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4739 OUT[5].t0 a_44640_1944.t23 VSS.t280 VSS.t279 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4740 VDD.t4231 a_26499_n2732 a_25895_n2624 VDD.t4230 pfet_06v0 ad=0.3975p pd=2.185u as=0.1521p ps=1.105u w=0.585u l=0.5u
X4741 VDD.t1069 a_21916_n6694.t21 a_30555_n2729 VDD.t1068 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X4742 a_46108_n2804 a_46020_n2760 VSS.t1271 VSS.t1270 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4743 a_11023_n4162.t10 a_13623_n4162.t45 VDD.t570 VDD.t569 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4744 VSS.t306 a_33496_n8222.t22 a_31548_n10172.t0 VSS.t305 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X4745 VSS.t898 a_4001_4292.t14 a_3935_4156.t2 VSS.t897 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X4746 a_29444_n4328.t5 a_29532_n4372.t9 VDD.t2055 VDD.t2054 pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
X4747 a_35804_n12212 a_35716_n12168 VSS.t2066 VSS.t2065 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4748 a_36140_n15781 a_36052_n15684 VSS.t4123 VSS.t4122 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4749 VDD.t1320 a_13623_n14874.t45 a_11023_n14874.t19 VDD.t1319 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4750 VDD.t2217 a_39724_n18917 a_39636_n18820 VDD.t2216 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4751 VDD.t538 a_23072_n13432.t101 a_25139_n2704 VDD.t537 pfet_06v0 ad=0.3432p pd=2.44u as=0.2028p ps=1.3u w=0.78u l=0.5u
X4752 a_38171_n3544 a_27225_n1572.t3 a_29263_n3588.t1 VSS.t3565 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X4753 a_32108_n2332.t8 a_35456_n4628.t22 VDD.t4095 VDD.t4094 pfet_06v0 ad=0.4392p pd=1.94u as=0.367p ps=1.92u w=1.22u l=0.5u
X4754 a_21692_n5468.t0 a_26440_n5940.t19 VSS.t365 VSS.t364 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X4755 VDD.t3456 a_35692_n17349 a_35604_n17252 VDD.t3455 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4756 a_45100_1467 a_45012_1564 VSS.t2640 VSS.t2639 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4757 VDD.t2469 a_32780_n18917 a_32692_n18820 VDD.t2468 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4758 VDD.t204 a_38256_1564.t23 OUT[3].t8 VDD.t203 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4759 VSS.t565 a_11023_n9518.t38 a_11087_n10138.t18 VSS.t64 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X4760 VDD.t3408 a_35692_n14213 a_35604_n14116 VDD.t2147 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4761 a_47116_n17349 a_47028_n17252 VSS.t3727 VSS.t3726 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4762 VDD.t3788 a_33452_n17349 a_33364_n17252 VDD.t3787 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4763 a_33900_n15348 a_33812_n15304 VSS.t4343 VSS.t4153 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4764 a_40196_1944 a_39748_2475 VDD.t1487 VDD.t1486 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X4765 a_37260_n7941 a_37172_n7844 VSS.t4144 VSS.t4143 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4766 a_11087_n10138.t19 a_11023_n9518.t39 VSS.t566 VSS.t66 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4767 VDD.t2488 a_28076_n18484 a_27988_n18440 VDD.t2487 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4768 VDD.t3245 a_27628_n3841 a_27540_n3797 VDD.t3244 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X4769 a_31961_n11340 a_23072_n13432.t102 VDD.t540 VDD.t539 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X4770 VDD.t3691 a_24569_n11820 a_24464_n11680 VDD.t3690 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X4771 VDD.t2473 a_30540_n18917 a_30452_n18820 VDD.t2472 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4772 a_41292_n17349 a_41204_n17252 VSS.t2234 VSS.t2233 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4773 a_47116_n14213 a_47028_n14116 VSS.t2236 VSS.t2235 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4774 VDD.t2728 a_33452_n14213 a_33364_n14116 VDD.t2727 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4775 a_21772_n452.t3 a_23564_n452.t9 VSS.t3749 VSS.t3748 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4776 a_40172_n17349 a_40084_n17252 VSS.t2287 VSS.t2286 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4777 a_41292_n14213 a_41204_n14116 VSS.t2259 VSS.t2258 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4778 a_31628_n5940.t16 a_33496_n6659.t39 VDD.t188 VDD.t187 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4779 VDD.t3938 a_31212_n17349 a_31124_n17252 VDD.t3937 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4780 a_13623_n22908.t3 a_21772_n452.t19 VDD.t1600 VDD.t1599 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4781 a_32085_n8248 a_31965_n8292 a_31341_n8292 VSS.t1629 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X4782 a_40172_n14213 a_40084_n14116 VSS.t1254 VSS.t1253 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4783 VDD.t60 a_45648_1564.t22 EOC.t8 VDD.t59 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4784 EOC.t0 a_45648_1564.t23 VSS.t43 VSS.t42 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4785 VDD.t2789 a_22588_n2020 a_22500_n1976 VDD.t2788 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4786 a_11087_n7460.t9 a_13623_n6840.t45 a_13501_n6460.t2 VSS.t746 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4787 a_13623_n17552.t8 a_21772_n8292.t23 VDD.t64 VDD.t63 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4788 a_27154_n9240 a_26470_n9322 VDD.t3131 VDD.t996 pfet_06v0 ad=61.199993f pd=0.7u as=0.1656p ps=1.28u w=0.36u l=0.5u
X4789 VDD.t2252 a_43644_n10644 a_43556_n10600 VDD.t2251 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4790 a_33920_n4 a_33820_n452.t3 VDD.t3802 VDD.t3801 pfet_06v0 ad=0.1464p pd=1.46u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4791 a_33608_n4284 a_33120_n3884 a_33868_n4240 VDD.t1079 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X4792 a_33776_n5896.t3 a_31628_n5940.t45 VDD.t154 VDD.t153 pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X4793 VSS.t4099 a_22968_n6679 a_22668_n14864.t0 VSS.t4098 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X4794 VDD.t3890 a_45660_n20052 a_45572_n20008 VDD.t3889 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4795 VDD.t385 a_10778_2852.t34 a_10712_4516.t20 VDD.t384 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X4796 a_29444_n4328.t2 a_29920_n3900.t22 VDD.t618 VDD.t617 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X4797 a_26981_n9010 a_26861_n8567 VDD.t2927 VDD.t2926 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X4798 VDD.t3008 a_44092_n9076 a_44004_n9032 VDD.t3007 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4799 VDD.t3280 a_41404_n10644 a_41316_n10600 VDD.t3279 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4800 VDD.t4296 a_44540_n20052 a_44452_n20008 VDD.t1293 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4801 VDD.t2037 a_43532_n7941 a_43444_n7844 VDD.t2036 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4802 VDD.t2710 a_43532_n4805 a_43444_n4708 VDD.t2709 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4803 VDD.t3928 a_42300_n20052 a_42212_n20008 VDD.t3927 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4804 a_28849_n13252 a_22220_690.t17 a_28645_n13252 VSS.t838 nfet_06v0 ad=0.1312p pd=1.14u as=0.1722p ps=1.24u w=0.82u l=0.6u
X4805 a_47197_908 a_43644_n705 VSS.t2842 VSS.t2841 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4806 a_26499_n2732 a_25795_n2716.t7 a_26915_n2672 VDD.t2358 pfet_06v0 ad=0.19315p pd=1.27u as=0.101p ps=0.905u w=0.505u l=0.5u
X4807 a_39948_n6373 a_39860_n6276 VSS.t2265 VSS.t2264 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4808 a_32560_n7020 a_31548_n10172.t25 VDD.t284 VDD.t283 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X4809 a_43644_n16916 a_43556_n16872 VSS.t1337 VSS.t1336 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4810 a_23072_n13432.t5 a_29744_n15604.t22 VDD.t1651 VDD.t1650 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X4811 VDD.t3530 a_40508_n4805 a_40420_n4708 VDD.t1455 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4812 a_24815_n3588.t0 a_29920_n3900.t23 VSS.t659 VSS.t658 nfet_06v0 ad=0.1248p pd=1u as=0.1248p ps=1u w=0.48u l=0.6u
X4813 VDD.t3617 a_34649_n2412 a_34544_n2272 VDD.t3616 pfet_06v0 ad=0.33755p pd=1.955u as=0.1313p ps=1.025u w=0.505u l=0.5u
X4814 a_11087_n23528.t61 a_2167_3472.t41 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X4815 VSS.t1937 a_24233_n3980 a_24128_n3840 VSS.t1936 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X4816 a_41404_n16916 a_41316_n16872 VSS.t1227 VSS.t1226 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4817 VDD.t2998 a_22588_n15781 a_22500_n15684 VDD.t2997 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4818 a_n263_3472.t8 a_22444_2253.t23 VDD.t2346 VDD.t2345 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4819 a_22444_332.t6 a_27259_804.t17 VDD.t812 VDD.t811 pfet_06v0 ad=0.52205p pd=2.045u as=0.30535p ps=1.605u w=0.985u l=0.5u
X4820 VSS.t709 a_29800_n5940.t22 a_28156_n6412.t0 VSS.t708 nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X4821 a_34176_n6976 a_32560_n7020 a_33048_n7420 VSS.t1330 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4822 a_29560_n3544 a_27259_804.t18 a_22444_332.t5 VSS.t858 nfet_06v0 ad=0.2132p pd=1.34u as=0.4161p ps=1.905u w=0.82u l=0.6u
X4823 VDD.t2456 a_28748_n18917 a_28660_n18820 VDD.t2455 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4824 a_34176_n3840 a_24481_761.t94 VSS.t830 VSS.t829 nfet_06v0 ad=43.199997f pd=0.6u as=0.2016p ps=1.48u w=0.36u l=0.6u
X4825 a_33572_n10980 a_28435_n10599 VDD.t3090 VDD.t3089 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X4826 VDD.t2401 a_23932_n16916 a_23844_n16872 VDD.t2400 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4827 VDD.t853 a_21772_n3588.t19 a_13623_n20230.t8 VDD.t852 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4828 VSS.t2659 a_21692_n5111.t5 a_21604_n5067 VSS.t404 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X4829 a_34372_n5112 a_24815_n3588.t23 a_34188_n5112 VSS.t27 nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X4830 VSS.t886 a_33776_n5896.t22 a_34708_n5896.t0 VSS.t885 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X4831 a_41292_n7941 a_41204_n7844 VSS.t3894 VSS.t3893 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4832 VDD.t2458 a_26508_n18917 a_26420_n18820 VDD.t2457 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4833 VDD.t435 a_33216_1944.t23 OUT[1].t8 VDD.t434 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4834 VDD.t1478 a_30808_n6334 a_30616_n6221 VDD.t1477 pfet_06v0 ad=0.2222p pd=1.89u as=0.2424p ps=1.465u w=0.505u l=0.5u
X4835 a_24180_n5112 a_24672_n11339 a_22220_n9860 VSS.t1966 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X4836 VDD.t3412 a_23564_1116.t9 a_21772_1116.t0 VDD.t2347 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X4837 a_30716_n1148 a_30408_n1104 VDD.t3653 VDD.t3652 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X4838 a_29444_n4328.t1 a_27259_804.t19 VDD.t814 VDD.t813 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X4839 a_23816_n10112 a_21604_n10116 a_22876_n10556 VDD.t3363 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X4840 VDD.t1805 a_44764_n1669 a_44676_n1572 VDD.t1804 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X4841 a_47116_n4805 a_47028_n4708 VSS.t2483 VSS.t2482 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X4842 VDD.t2437 a_26531_n10207 a_26239_n11428 VDD.t2436 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X4843 VSS.t642 a_13623_n20230.t45 a_11023_n20230.t0 VSS.t641 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
D135 VSS.t367 a_26388_n17606.t13 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X4844 a_27205_n16088 a_27085_n16132 VSS.t1957 VSS.t1956 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X4845 a_35916_n4 a_35816_n174 VDD.t3308 VDD.t3307 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X4846 VSS.t554 a_23072_n13432.t103 a_23024_n704 VSS.t553 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
R0 VDD.t2117 VDD.t529 593.75
R1 VDD.t4046 VDD.t506 570.602
R2 VDD.t3443 VDD.t1953 527.779
R3 VDD.t2657 VDD.n1339 525.553
R4 VDD.t3400 VDD.t2023 518.519
R5 VDD.t1502 VDD.t2657 518.519
R6 VDD.t2440 VDD.t1502 518.519
R7 VDD.t1158 VDD.t2440 518.519
R8 VDD.t2194 VDD.t1158 518.519
R9 VDD.t3037 VDD.t2194 518.519
R10 VDD.t2548 VDD.t3037 518.519
R11 VDD.t3068 VDD.t1804 518.519
R12 VDD.t3295 VDD.t3068 518.519
R13 VDD.t3320 VDD.t2307 518.519
R14 VDD.t3614 VDD.t1455 518.519
R15 VDD.t1455 VDD.t1546 518.519
R16 VDD.t1546 VDD.t2228 518.519
R17 VDD.t2228 VDD.t2794 518.519
R18 VDD.t3098 VDD.t3001 518.519
R19 VDD.t2677 VDD.t4181 518.519
R20 VDD.t2707 VDD.t3043 518.519
R21 VDD.t2323 VDD.t3626 518.519
R22 VDD.t2266 VDD.t2323 518.519
R23 VDD.t2147 VDD.t2266 518.519
R24 VDD.t1368 VDD.t2147 518.519
R25 VDD.t1419 VDD.t1368 518.519
R26 VDD.t1218 VDD.t2997 518.519
R27 VDD.t1787 VDD.t1218 518.519
R28 VDD.t3644 VDD.t988 518.519
R29 VDD.t988 VDD.t2776 518.519
R30 VDD.t2776 VDD.t2366 518.519
R31 VDD.t2366 VDD.t953 518.519
R32 VDD.t953 VDD.t1201 518.519
R33 VDD.t1201 VDD.t1328 518.519
R34 VDD.t1328 VDD.t2385 518.519
R35 VDD.t2385 VDD.t3144 518.519
R36 VDD.t931 VDD.t914 518.519
R37 VDD.t2233 VDD.t3716 518.519
R38 VDD.t2455 VDD.t2510 518.519
R39 VDD.t1584 VDD.t3538 518.519
R40 VDD.t1607 VDD.t1584 518.519
R41 VDD.t3554 VDD.t1607 518.519
R42 VDD.t3335 VDD.t3554 518.519
R43 VDD.t3343 VDD.t3335 518.519
R44 VDD.t1239 VDD.t3343 518.519
R45 VDD.t1609 VDD.t1239 518.519
R46 VDD.t908 VDD.t1609 518.519
R47 VDD.t3563 VDD.t2044 518.519
R48 VDD.t2044 VDD.t986 518.519
R49 VDD.t986 VDD.t2192 518.519
R50 VDD.t2192 VDD.t3011 518.519
R51 VDD.t3011 VDD.t961 518.519
R52 VDD.t961 VDD.t2778 518.519
R53 VDD.t2094 VDD.t1002 518.519
R54 VDD.t1002 VDD.t1461 518.519
R55 VDD.t1461 VDD.t2086 518.519
R56 VDD.t2086 VDD.t2218 518.519
R57 VDD.t2218 VDD.t2792 518.519
R58 VDD.t2792 VDD.t1162 518.519
R59 VDD.t1162 VDD.t2048 518.519
R60 VDD.t3351 VDD.t4055 518.519
R61 VDD.t641 VDD.t4057 515.047
R62 VDD.t2956 VDD.t2260 510.418
R63 VDD.t1947 VDD.t1734 506.945
R64 VDD.t1398 VDD.t1157 504.63
R65 VDD.t3256 VDD.t394 497.685
R66 VDD.t349 VDD.t4112 496.529
R67 VDD.t1082 VDD.t633 493.057
R68 VDD.t519 VDD.t3026 488.426
R69 VDD.n269 VDD.t2968 483.796
R70 VDD.t281 VDD.t4139 483.796
R71 VDD.t1446 VDD.t743 478.01
R72 VDD.t3275 VDD.t4257 474.538
R73 VDD.n517 VDD.t4 472.223
R74 VDD.t3795 VDD.t3911 472.223
R75 VDD.t2393 VDD.t480 472.223
R76 VDD.t2295 VDD.t4064 472.223
R77 VDD.t2733 VDD.t2442 468.75
R78 VDD.t1395 VDD.t2319 460.649
R79 VDD.t4033 VDD.t2993 460.649
R80 VDD.n534 VDD.t1594 453.786
R81 VDD.n1670 VDD.t858 453.786
R82 VDD.t2168 VDD.t1269 453.704
R83 VDD.t1927 VDD.t155 453.704
R84 VDD.t2438 VDD.t710 451.389
R85 VDD.n510 VDD.t3053 447.918
R86 VDD.t529 VDD.t3766 440.973
R87 VDD.t753 VDD.t137 437.5
R88 VDD.t2794 VDD.t324 435.185
R89 VDD.t3610 VDD.t703 435.185
R90 VDD.t4118 VDD.t2636 435.185
R91 VDD.t4117 VDD.t2370 435.185
R92 VDD.t4060 VDD.t2753 435.185
R93 VDD.t3204 VDD.t3 435.185
R94 VDD.t1132 VDD.t522 435.185
R95 VDD.t496 VDD.t1419 435.185
R96 VDD.t2457 VDD.t4062 435.185
R97 VDD.n2024 VDD.t3638 430.623
R98 VDD.t3650 VDD.t530 429.399
R99 VDD.t2416 VDD.t2622 425.926
R100 VDD.t1853 VDD.t2103 422.454
R101 VDD.t1151 VDD.t3608 421.296
R102 VDD.t3580 VDD.t1082 416.668
R103 VDD.t634 VDD.t472 415.51
R104 VDD.t443 VDD.t4121 414.353
R105 VDD.t467 VDD.t2932 406.587
R106 VDD.t804 VDD.t3234 403.935
R107 VDD.t3760 VDD.t2592 403.935
R108 VDD.t2189 VDD.t1548 402.779
R109 VDD.t1622 VDD.t2503 402.779
R110 VDD.t2033 VDD.t3309 402.779
R111 VDD.n2116 VDD.t1787 396.068
R112 VDD.n223 VDD.t908 396.068
R113 VDD.n2175 VDD.t1662 395.916
R114 VDD.n2287 VDD.t3774 395.916
R115 VDD.t2023 VDD.n1385 395.841
R116 VDD.t4294 VDD.n1261 395.841
R117 VDD.t2249 VDD.n1220 395.841
R118 VDD.t4290 VDD.n1174 395.841
R119 VDD.t2522 VDD.n1088 395.841
R120 VDD.t4282 VDD.n1041 395.841
R121 VDD.t2798 VDD.n994 395.841
R122 VDD.t3419 VDD.n914 395.841
R123 VDD.t3049 VDD.n867 395.841
R124 VDD.t2007 VDD.n820 395.841
R125 VDD.t3449 VDD.n741 395.841
R126 VDD.t2864 VDD.n694 395.841
R127 VDD.t3544 VDD.t2663 388.889
R128 VDD.n1386 VDD.t3770 388.889
R129 VDD.n1340 VDD.t2548 388.889
R130 VDD.t3206 VDD.t2759 388.889
R131 VDD.t3045 VDD.t3578 388.889
R132 VDD.t3836 VDD.t2780 388.889
R133 VDD.t3464 VDD.t982 388.889
R134 VDD.t1580 VDD.t1214 388.889
R135 VDD.t2681 VDD.t2025 388.889
R136 VDD.t2307 VDD.t4288 388.889
R137 VDD.t3333 VDD.t2817 388.889
R138 VDD.t2149 VDD.t2569 388.889
R139 VDD.t1887 VDD.t2782 388.889
R140 VDD.t3513 VDD.t2481 388.889
R141 VDD.t2890 VDD.t2679 388.889
R142 VDD.t3085 VDD.t1435 388.889
R143 VDD.t941 VDD.t3303 388.889
R144 VDD.t3316 VDD.t2755 388.889
R145 VDD.t2182 VDD.t2151 388.889
R146 VDD.t2391 VDD.t3747 388.889
R147 VDD.t2134 VDD.t2129 388.889
R148 VDD.t2888 VDD.t2363 388.889
R149 VDD.t1986 VDD.t3821 388.889
R150 VDD.t3202 VDD.t3915 388.889
R151 VDD.t893 VDD.t3846 388.889
R152 VDD.t3531 VDD.t893 388.889
R153 VDD.t3417 VDD.t1500 388.889
R154 VDD.t3873 VDD.t957 388.889
R155 VDD.t3913 VDD.t2709 388.889
R156 VDD.t2673 VDD.t3793 388.889
R157 VDD.t2071 VDD.t2539 388.889
R158 VDD.t1537 VDD.t1431 388.889
R159 VDD.t1116 VDD.t2934 388.889
R160 VDD.t3614 VDD.t2558 388.889
R161 VDD.t3173 VDD.t3789 388.889
R162 VDD.t3246 VDD.t4211 388.889
R163 VDD.t1354 VDD.t1473 388.889
R164 VDD.t2013 VDD.t4266 388.889
R165 VDD.t2483 VDD.t1207 388.889
R166 VDD.t2395 VDD.t3250 388.889
R167 VDD.t3001 VDD.t3132 388.889
R168 VDD.n1175 VDD.t969 388.889
R169 VDD.t2291 VDD.t1626 388.889
R170 VDD.t2380 VDD.t2912 388.889
R171 VDD.t3341 VDD.t2031 388.889
R172 VDD.t3117 VDD.t1912 388.889
R173 VDD.t3453 VDD.t1922 388.889
R174 VDD.t1411 VDD.t3939 388.889
R175 VDD.t967 VDD.t1722 388.889
R176 VDD.t2898 VDD.t967 388.889
R177 VDD.t4020 VDD.t1443 388.889
R178 VDD.t1992 VDD.t1857 388.889
R179 VDD.t1339 VDD.t2036 388.889
R180 VDD.t2321 VDD.t4183 388.889
R181 VDD.t2942 VDD.t4105 388.889
R182 VDD.t3398 VDD.t4053 388.889
R183 VDD.t3070 VDD.t1840 388.889
R184 VDD.t4181 VDD.t3811 388.889
R185 VDD.t3524 VDD.t2665 388.889
R186 VDD.t3967 VDD.t2790 388.889
R187 VDD.t3129 VDD.t2874 388.889
R188 VDD.t2444 VDD.t4072 388.889
R189 VDD.t1523 VDD.t1358 388.889
R190 VDD.t3406 VDD.t2269 388.889
R191 VDD.t2112 VDD.t1235 388.889
R192 VDD.t3799 VDD.t3803 388.889
R193 VDD.t1914 VDD.t2119 388.889
R194 VDD.t4276 VDD.t2027 388.889
R195 VDD.t998 VDD.t3248 388.889
R196 VDD.t3567 VDD.t2868 388.889
R197 VDD.t4040 VDD.t1291 388.889
R198 VDD.t2583 VDD.t3576 388.889
R199 VDD.t2330 VDD.t2583 388.889
R200 VDD.t3007 VDD.t1865 388.889
R201 VDD.t3682 VDD.t2675 388.889
R202 VDD.t3108 VDD.t3154 388.889
R203 VDD.t975 VDD.t3515 388.889
R204 VDD.t2359 VDD.t3353 388.889
R205 VDD.t3142 VDD.t1409 388.889
R206 VDD.t4068 VDD.t2659 388.889
R207 VDD.t1130 VDD.t3751 388.889
R208 VDD.t1130 VDD.t2127 388.889
R209 VDD.t3522 VDD.t2546 388.889
R210 VDD.t2299 VDD.t3634 388.889
R211 VDD.t3853 VDD.t3262 388.889
R212 VDD.t1415 VDD.t3885 388.889
R213 VDD.t1910 VDD.t4197 388.889
R214 VDD.t1233 VDD.t3384 388.889
R215 VDD.t2590 VDD.t2809 388.889
R216 VDD.t3311 VDD.t2370 388.889
R217 VDD.t1789 VDD.t3745 388.889
R218 VDD.t2729 VDD.t2962 388.889
R219 VDD.t2896 VDD.t2870 388.889
R220 VDD.t2214 VDD.t1510 388.889
R221 VDD.t2667 VDD.t2038 388.889
R222 VDD.t977 VDD.t3893 388.889
R223 VDD.t2774 VDD.t1628 388.889
R224 VDD.t4038 VDD.t2774 388.889
R225 VDD.t2368 VDD.t3198 388.889
R226 VDD.t2251 VDD.t2361 388.889
R227 VDD.t2253 VDD.t2669 388.889
R228 VDD.t1682 VDD.t3949 388.889
R229 VDD.t2860 VDD.t4042 388.889
R230 VDD.t1231 VDD.t4096 388.889
R231 VDD.t3279 VDD.t2489 388.889
R232 VDD.t1439 VDD.t3686 388.889
R233 VDD.t1439 VDD.t2493 388.889
R234 VDD.t1800 VDD.t2757 388.889
R235 VDD.t3574 VDD.t3572 388.889
R236 VDD.t1812 VDD.t4199 388.889
R237 VDD.t2101 VDD.t2277 388.889
R238 VDD.t3087 VDD.t2450 388.889
R239 VDD.t3986 VDD.t1718 388.889
R240 VDD.t2807 VDD.t3586 388.889
R241 VDD.t1810 VDD.t3204 388.889
R242 VDD.t4207 VDD.t3591 388.889
R243 VDD.t1481 VDD.t1134 388.889
R244 VDD.t2800 VDD.t3074 388.889
R245 VDD.t4201 VDD.t1582 388.889
R246 VDD.t898 VDD.t1138 388.889
R247 VDD.t4213 VDD.t2725 388.889
R248 VDD.t2940 VDD.t3081 388.889
R249 VDD.t3941 VDD.t2940 388.889
R250 VDD.t3318 VDD.t1620 388.889
R251 VDD.t2843 VDD.t3947 388.889
R252 VDD.t1212 VDD.t2420 388.889
R253 VDD.t3988 VDD.t1423 388.889
R254 VDD.t1707 VDD.t1535 388.889
R255 VDD.t3838 VDD.t1937 388.889
R256 VDD.t3238 VDD.t3162 388.889
R257 VDD.t3043 VDD.t2092 388.889
R258 VDD.t4238 VDD.t2201 388.889
R259 VDD.t2823 VDD.t3832 388.889
R260 VDD.t2301 VDD.t1889 388.889
R261 VDD.t3187 VDD.t3421 388.889
R262 VDD.t3290 VDD.t2084 388.889
R263 VDD.t1730 VDD.t4232 388.889
R264 VDD.t2835 VDD.t984 388.889
R265 VDD.t2061 VDD.t2029 388.889
R266 VDD.t1777 VDD.t3369 388.889
R267 VDD.t1479 VDD.t1984 388.889
R268 VDD.t3015 VDD.t2554 388.889
R269 VDD.t3469 VDD.t1739 388.889
R270 VDD.t2157 VDD.t3640 388.889
R271 VDD.t4177 VDD.t3923 388.889
R272 VDD.t4171 VDD.t1259 388.889
R273 VDD.t1226 VDD.t2560 388.889
R274 VDD.t3112 VDD.t3665 388.889
R275 VDD.t2315 VDD.t4227 388.889
R276 VDD.t2125 VDD.t2315 388.889
R277 VDD.t3381 VDD.t4167 388.889
R278 VDD.t3688 VDD.t1245 388.889
R279 VDD.t3536 VDD.t1228 388.889
R280 VDD.t2721 VDD.t4011 388.889
R281 VDD.t3451 VDD.t2642 388.889
R282 VDD.t3345 VDD.t1297 388.889
R283 VDD.t3091 VDD.t1251 388.889
R284 VDD.t2526 VDD.t2172 388.889
R285 VDD.t2526 VDD.t1370 388.889
R286 VDD.t1679 VDD.t1195 388.889
R287 VDD.t3976 VDD.t939 388.889
R288 VDD.t965 VDD.t3528 388.889
R289 VDD.t3929 VDD.t3377 388.889
R290 VDD.t3999 VDD.t3252 388.889
R291 VDD.t1732 VDD.t2640 388.889
R292 VDD.t1737 VDD.t2520 388.889
R293 VDD.t3136 VDD.t3626 388.889
R294 VDD.t2209 VDD.t2829 388.889
R295 VDD.t2159 VDD.t2661 388.889
R296 VDD.t4280 VDD.t4286 388.889
R297 VDD.t1099 VDD.t2902 388.889
R298 VDD.t4076 VDD.t3102 388.889
R299 VDD.t2448 VDD.t2398 388.889
R300 VDD.t3156 VDD.t2303 388.889
R301 VDD.t3236 VDD.t3156 388.889
R302 VDD.t1632 VDD.t3881 388.889
R303 VDD.t1684 VDD.t2839 388.889
R304 VDD.t3842 VDD.t4101 388.889
R305 VDD.t3003 VDD.t1982 388.889
R306 VDD.t3277 VDD.t2954 388.889
R307 VDD.t1802 VDD.t1350 388.889
R308 VDD.t2900 VDD.t3005 388.889
R309 VDD.t3783 VDD.t3425 388.889
R310 VDD.t3783 VDD.t3152 388.889
R311 VDD.t2476 VDD.t1990 388.889
R312 VDD.t4218 VDD.t2042 388.889
R313 VDD.t3654 VDD.t4169 388.889
R314 VDD.t3718 VDD.t971 388.889
R315 VDD.t2402 VDD.t3477 388.889
R316 VDD.t2462 VDD.t4292 388.889
R317 VDD.t3013 VDD.t4158 388.889
R318 VDD.t1190 VDD.t3644 388.889
R319 VDD.n2103 VDD.t3144 388.889
R320 VDD.t3805 VDD.t3423 388.889
R321 VDD.t3642 VDD.t1332 388.889
R322 VDD.t4163 VDD.t3963 388.889
R323 VDD.t4156 VDD.t1616 388.889
R324 VDD.t1224 VDD.t3995 388.889
R325 VDD.t3110 VDD.t3041 388.889
R326 VDD.t2255 VDD.t4225 388.889
R327 VDD.t2275 VDD.t2255 388.889
R328 VDD.t1761 VDD.t4150 388.889
R329 VDD.t1289 VDD.t1097 388.889
R330 VDD.t2944 VDD.t1417 388.889
R331 VDD.t2297 VDD.t1832 388.889
R332 VDD.t3178 VDD.t2372 388.889
R333 VDD.t3636 VDD.t933 388.889
R334 VDD.t1179 VDD.t1247 388.889
R335 VDD.t4272 VDD.t2063 388.889
R336 VDD.t1249 VDD.t4272 388.889
R337 VDD.t2207 VDD.t2652 388.889
R338 VDD.t1388 VDD.t1421 388.889
R339 VDD.t1674 VDD.t2485 388.889
R340 VDD.t3373 VDD.t2991 388.889
R341 VDD.t2703 VDD.t3971 388.889
R342 VDD.t2603 VDD.t1724 388.889
R343 VDD.t2422 VDD.t3427 388.889
R344 VDD.t1785 VDD.t2872 388.889
R345 VDD.t4103 VDD.t1785 388.889
R346 VDD.t3158 VDD.t2533 388.889
R347 VDD.t3671 VDD.t1975 388.889
R348 VDD.t2575 VDD.t3455 388.889
R349 VDD.t3435 VDD.t1433 388.889
R350 VDD.t3266 VDD.t3404 388.889
R351 VDD.t3584 VDD.t2537 388.889
R352 VDD.t3034 VDD.t3484 388.889
R353 VDD.t931 VDD.t3787 388.889
R354 VDD.t1241 VDD.t3240 388.889
R355 VDD.t3809 VDD.t2815 388.889
R356 VDD.t923 VDD.t3100 388.889
R357 VDD.t3937 VDD.t4203 388.889
R358 VDD.t3379 VDD.t959 388.889
R359 VDD.t1345 VDD.t1471 388.889
R360 VDD.t1900 VDD.t4270 388.889
R361 VDD.t4005 VDD.t2831 388.889
R362 VDD.t3673 VDD.t1557 388.889
R363 VDD.t2821 VDD.t3119 388.889
R364 VDD.t1321 VDD.t3371 388.889
R365 VDD.t3708 VDD.t1186 388.889
R366 VDD.t3867 VDD.t3708 388.889
R367 VDD.t2958 VDD.t2849 388.889
R368 VDD.t918 VDD.t2414 388.889
R369 VDD.t927 VDD.t3712 388.889
R370 VDD.t2979 VDD.t935 388.889
R371 VDD.t1343 VDD.t1498 388.889
R372 VDD.t2579 VDD.t3441 388.889
R373 VDD.t3917 VDD.t3593 388.889
R374 VDD.t3439 VDD.t1136 388.889
R375 VDD.t3439 VDD.t1979 388.889
R376 VDD.t2404 VDD.t1539 388.889
R377 VDD.t2833 VDD.t2216 388.889
R378 VDD.t2966 VDD.t3160 388.889
R379 VDD.t4143 VDD.t2845 388.889
R380 VDD.t1149 VDD.t3164 388.889
R381 VDD.t3367 VDD.t1437 388.889
R382 VDD.t2491 VDD.t1793 388.889
R383 VDD.t3935 VDD.t2811 388.889
R384 VDD.t2894 VDD.t2811 388.889
R385 VDD.t3827 VDD.t3830 388.889
R386 VDD.t1945 VDD.t3305 388.889
R387 VDD.t1634 VDD.t904 388.889
R388 VDD.t3166 VDD.t3778 388.889
R389 VDD.t1898 VDD.t3877 388.889
R390 VDD.t1280 VDD.t874 388.889
R391 VDD.t1103 VDD.t3171 388.889
R392 VDD.t3943 VDD.t2516 388.889
R393 VDD.t2468 VDD.t3943 388.889
R394 VDD.t1105 VDD.t2271 388.889
R395 VDD.t3314 VDD.t2203 388.889
R396 VDD.t3180 VDD.t2153 388.889
R397 VDD.t1575 VDD.t2090 388.889
R398 VDD.t2472 VDD.t2220 388.889
R399 VDD.t3169 VDD.t2273 388.889
R400 VDD.t3146 VDD.t2264 388.889
R401 VDD.t2510 VDD.t2571 388.889
R402 VDD.t1142 VDD.t2457 388.889
R403 VDD.t2174 VDD.t1988 388.889
R404 VDD.t3538 VDD.t1969 388.889
R405 VDD.t1293 VDD.n651 388.889
R406 VDD.n652 VDD.t1293 388.889
R407 VDD.n653 VDD.t3563 388.889
R408 VDD.t2778 VDD.n219 388.889
R409 VDD.n218 VDD.t2094 388.889
R410 VDD.n2277 VDD.t2048 388.889
R411 VDD.t1341 VDD.t4001 388.889
R412 VDD.t2585 VDD.n2281 388.889
R413 VDD.t1916 VDD.t651 384.26
R414 VDD.t2886 VDD.t2452 381.945
R415 VDD.t980 VDD.t2928 381.945
R416 VDD.t3973 VDD.t880 381.945
R417 VDD.t3077 VDD.t3534 381.945
R418 VDD.t3297 VDD.t2161 380.788
R419 VDD.n1097 VDD.t1197 379.075
R420 VDD.n2114 VDD.t937 379.075
R421 VDD.t912 VDD.t2731 373.844
R422 VDD.t973 VDD.t1779 373.022
R423 VDD.t1517 VDD.t4154 371.529
R424 VDD.t1774 VDD.t1475 370.37
R425 VDD.t2784 VDD.t747 365.741
R426 VDD.t1459 VDD.t773 365.741
R427 VDD.t3182 VDD.t473 365.741
R428 VDD.t2556 VDD.t461 365.741
R429 VDD.t3772 VDD.t483 365.741
R430 VDD.t3242 VDD.t1025 364.92
R431 VDD.t2231 VDD.t1977 364.92
R432 VDD.t3595 VDD.t1092 363.426
R433 VDD.n566 VDD.t3375 362.269
R434 VDD.n576 VDD.t1253 362.269
R435 VDD.n1776 VDD.t2906 362.269
R436 VDD.n1612 VDD.t358 361.286
R437 VDD.n447 VDD.t398 361.286
R438 VDD.n1509 VDD.t3768 361.192
R439 VDD.n1967 VDD.t2630 361.192
R440 VDD.n279 VDD.t2628 361.192
R441 VDD.n351 VDD.t2632 361.178
R442 VDD.n1795 VDD.t364 361.132
R443 VDD.t2065 VDD.t1027 361.111
R444 VDD.n525 VDD.t3349 358.76
R445 VDD.t1489 VDD.t4044 355.437
R446 VDD.t2188 VDD.t1 355.437
R447 VDD.t396 VDD.n560 354.168
R448 VDD.n1598 VDD.t360 354.168
R449 VDD.n1604 VDD.t796 354.168
R450 VDD.t4240 VDD.t3212 351.853
R451 VDD.t1449 VDD.t746 350.695
R452 VDD.t1365 VDD.t2910 348.865
R453 VDD.t1971 VDD.t2786 348.865
R454 VDD.t4030 VDD.t3473 348.865
R455 VDD.t2989 VDD.t1504 348.865
R456 VDD.t4141 VDD.t527 347.223
R457 VDD.t173 VDD.t611 347.223
R458 VDD.t1508 VDD.t2862 346.065
R459 VDD.t503 VDD.t2825 346.065
R460 VDD.n586 VDD.t2430 344.908
R461 VDD.t2841 VDD.t3519 344.908
R462 VDD.t2211 VDD.t2040 344.908
R463 VDD.t794 VDD.t2981 342.892
R464 VDD.t718 VDD.t2719 342.594
R465 VDD.t642 VDD.t1769 342.594
R466 VDD.t1265 VDD.t3558 342.594
R467 VDD.t1495 VDD.t3652 341.772
R468 VDD.t2459 VDD.t490 340.279
R469 VDD.t2825 VDD.t2244 340.279
R470 VDD.t805 VDD.n1265 339.12
R471 VDD.n2104 VDD.t3598 339.12
R472 VDD.n1858 VDD.t4274 337.969
R473 VDD.t963 VDD.t2436 337.964
R474 VDD.t3057 VDD.n601 331.019
R475 VDD.t1850 VDD.t4220 331.019
R476 VDD.t2389 VDD.t3116 331.019
R477 VDD.t2313 VDD.t3076 331.019
R478 VDD.t3200 VDD.t2464 331.019
R479 VDD.t1483 VDD.t4028 329.861
R480 VDD.t2078 VDD.t1577 329.041
R481 VDD.t1101 VDD.t943 326.762
R482 VDD.t1040 VDD.t1048 326.264
R483 VDD.t2984 VDD.t418 325.231
R484 VDD.n139 VDD.t436 321.339
R485 VDD.n174 VDD.t843 321.065
R486 VDD.n116 VDD.t376 318.656
R487 VDD.t2550 VDD.t2082 318.399
R488 VDD.t2727 VDD.t1726 317.13
R489 VDD.n178 VDD.t339 316.43
R490 VDD.t3980 VDD.t1571 315.973
R491 VDD.n1669 VDD.t3892 315.853
R492 VDD.n919 VDD.t2857 314.815
R493 VDD.n7 VDD.t213 312.738
R494 VDD.n20 VDD.t1846 312.738
R495 VDD.n32 VDD.t2692 312.738
R496 VDD.n43 VDD.t115 312.738
R497 VDD.n55 VDD.t545 312.738
R498 VDD.n67 VDD.t130 312.738
R499 VDD.n79 VDD.t76 312.738
R500 VDD.n91 VDD.t401 312.738
R501 VDD.t1550 VDD.t3975 312.5
R502 VDD.t798 VDD.t756 312.353
R503 VDD.t3844 VDD.t3021 311.344
R504 VDD.n133 VDD.t2351 311.322
R505 VDD.n132 VDD.t2021 311.322
R506 VDD.n142 VDD.t2009 311.204
R507 VDD.n143 VDD.t2011 311.204
R508 VDD.n6 VDD.t226 311.132
R509 VDD.n19 VDD.t587 311.132
R510 VDD.n31 VDD.t561 311.132
R511 VDD.n42 VDD.t673 311.132
R512 VDD.n54 VDD.t269 311.132
R513 VDD.n66 VDD.t1743 311.132
R514 VDD.n78 VDD.t1317 311.132
R515 VDD.n90 VDD.t103 311.132
R516 VDD.t732 VDD.n502 309.14
R517 VDD.t4 VDD.t3028 307.87
R518 VDD.t1703 VDD.t738 307.87
R519 VDD.n1346 VDD.t11 305.557
R520 VDD.t19 VDD.t3520 305.557
R521 VDD.t3520 VDD.t643 305.557
R522 VDD.t3269 VDD.t777 305.557
R523 VDD.t3148 VDD.t3700 305.557
R524 VDD.t2530 VDD.t3677 303.241
R525 VDD.n1097 VDD.t848 301.887
R526 VDD.t236 VDD.t3753 300.926
R527 VDD.t4193 VDD.t3125 300.926
R528 VDD.n1857 VDD.t3192 299.769
R529 VDD.t780 VDD.t811 299.166
R530 VDD.t3504 VDD.t1605 296.296
R531 VDD.t2595 VDD.t2530 296.296
R532 VDD.t3990 VDD.t2478 294.505
R533 VDD.t2750 VDD.t1268 292.825
R534 VDD.t784 VDD.t479 292.825
R535 VDD.t1998 VDD.t2165 292.825
R536 VDD.t2544 VDD.t4111 292.825
R537 VDD.t2717 VDD.t3431 290.51
R538 VDD.t1124 VDD.t3602 290.51
R539 VDD.t43 VDD.t3961 290.51
R540 VDD.t695 VDD.t661 288.568
R541 VDD.t736 VDD.t3413 287.038
R542 VDD.t741 VDD.t3347 287.038
R543 VDD.t3540 VDD.t515 287.038
R544 VDD.t1660 VDD.t3462 287.038
R545 VDD.t1031 VDD.t1237 287.038
R546 VDD.t1153 VDD.t759 287.038
R547 VDD.t2950 VDD.t520 287.038
R548 VDD.t994 VDD.t501 287.038
R549 VDD.t4152 VDD.t2474 287.038
R550 VDD.t1569 VDD.t469 287.038
R551 VDD.t511 VDD.t1624 287.038
R552 VDD.t2683 VDD.t525 287.038
R553 VDD.t61 VDD.t1906 286.055
R554 VDD.t317 VDD.t1029 284.723
R555 VDD.t4059 VDD.t1519 283.565
R556 VDD.t1429 VDD.t1072 282.558
R557 VDD.t3287 VDD.t1941 282.408
R558 VDD.t2262 VDD.t3797 282.408
R559 VDD.t4084 VDD.t4088 282.408
R560 VDD.t4080 VDD.t4082 282.408
R561 VDD.t4094 VDD.t4090 282.408
R562 VDD.t293 VDD.t291 282.408
R563 VDD.t3638 VDD.t3486 282.408
R564 VDD.t2285 VDD.t2282 282.408
R565 VDD.t1646 VDD.t1648 282.408
R566 VDD.t1650 VDD.t1638 282.408
R567 VDD.t1636 VDD.t1642 282.408
R568 VDD.t715 VDD.t761 282.408
R569 VDD.t1885 VDD.t2851 281.25
R570 VDD.t4234 VDD.t2358 280.094
R571 VDD.t3232 VDD.t2241 278.115
R572 VDD.t1107 VDD.t3834 277.779
R573 VDD.t2764 VDD.t1330 277.779
R574 VDD.t2410 VDD.t3079 277.779
R575 VDD.t1282 VDD.t3327 277.779
R576 VDD.t1613 VDD.t4230 277.779
R577 VDD.t1475 VDD.t1796 277.779
R578 VDD.t1465 VDD.t3499 277.779
R579 VDD.t2099 VDD.t2599 277.779
R580 VDD.t3701 VDD.t2877 277.779
R581 VDD.n2174 VDD.t2599 275.464
R582 VDD.t1765 VDD.t3694 273.149
R583 VDD.t1798 VDD.t139 273.149
R584 VDD.t507 VDD.t1676 273.149
R585 VDD.t3933 VDD.t3259 271.991
R586 VDD.t3194 VDD.t844 271.991
R587 VDD.t1081 VDD.t792 270.834
R588 VDD.t1796 VDD.t3985 270.834
R589 VDD.n1949 VDD.t4179 270.012
R590 VDD.t713 VDD.t2397 268.519
R591 VDD.t481 VDD.t689 268.519
R592 VDD.t3899 VDD.t3905 267.623
R593 VDD.t1177 VDD.t1175 267.623
R594 VDD.t1666 VDD.t1668 267.623
R595 VDD.t3739 VDD.t3737 267.623
R596 VDD.t4262 VDD.t1544 267.361
R597 VDD.n325 VDD.t1118 267.361
R598 VDD.t1935 VDD.t1287 267.361
R599 VDD.t3482 VDD.t1164 266.985
R600 VDD.t3628 VDD.n1508 266.204
R601 VDD.n1098 VDD.t751 266.204
R602 VDD.t925 VDD.t3264 265.83
R603 VDD.t3460 VDD.t2946 265.046
R604 VDD.n441 VDD.t2246 265.046
R605 VDD.t2178 VDD.t846 265.046
R606 VDD.t2910 VDD.t3667 261.911
R607 VDD.t890 VDD.t1705 259.26
R608 VDD.t2349 VDD.t2334 259.26
R609 VDD.t2347 VDD.t2349 259.26
R610 VDD.t2343 VDD.t2347 259.26
R611 VDD.t2345 VDD.t2343 259.26
R612 VDD.t2340 VDD.t2345 259.26
R613 VDD.t457 VDD.t2340 259.26
R614 VDD.t459 VDD.t457 259.26
R615 VDD.t451 VDD.t459 259.26
R616 VDD.t453 VDD.t451 259.26
R617 VDD.t455 VDD.t453 259.26
R618 VDD.t619 VDD.t455 259.26
R619 VDD.t447 VDD.t619 259.26
R620 VDD.t3897 VDD.t3903 259.26
R621 VDD.t2711 VDD.t2715 259.26
R622 VDD.t1126 VDD.t1122 259.26
R623 VDD.t57 VDD.t45 259.26
R624 VDD.t45 VDD.t53 259.26
R625 VDD.t55 VDD.t49 259.26
R626 VDD.t239 VDD.t2495 259.26
R627 VDD.t2501 VDD.t2499 259.26
R628 VDD.t3059 VDD.t1781 259.26
R629 VDD.t199 VDD.t203 259.26
R630 VDD.t193 VDD.t197 259.26
R631 VDD.t1694 VDD.t1686 259.26
R632 VDD.t1654 VDD.t1658 259.26
R633 VDD.t1658 VDD.t1652 259.26
R634 VDD.t1599 VDD.t1592 259.26
R635 VDD.t1588 VDD.t1597 259.26
R636 VDD.t1590 VDD.t779 259.26
R637 VDD.t1390 VDD.t1392 259.26
R638 VDD.t2650 VDD.t2766 259.26
R639 VDD.t1270 VDD.t2987 259.26
R640 VDD.t782 VDD.t12 259.26
R641 VDD.t738 VDD.t782 259.26
R642 VDD.t4131 VDD.t1703 259.26
R643 VDD.t2803 VDD.t2805 259.26
R644 VDD.t876 VDD.t3511 259.26
R645 VDD.t2916 VDD.t2918 259.26
R646 VDD.t856 VDD.t575 259.26
R647 VDD.t850 VDD.t571 259.26
R648 VDD.t1046 VDD.t3024 259.26
R649 VDD.t1070 VDD.t3727 259.26
R650 VDD.t3733 VDD.t3729 259.26
R651 VDD.n1262 VDD.t1020 259.26
R652 VDD.t2755 VDD.n1262 259.26
R653 VDD.t3698 VDD.t3551 259.26
R654 VDD.t3494 VDD.t4065 259.26
R655 VDD.t3969 VDD.t3098 259.26
R656 VDD.t3883 VDD.t3969 259.26
R657 VDD.t3556 VDD.t3883 259.26
R658 VDD.t2446 VDD.t3556 259.26
R659 VDD.t3549 VDD.t2446 259.26
R660 VDD.t3134 VDD.t3549 259.26
R661 VDD.t1630 VDD.t3134 259.26
R662 VDD.t2418 VDD.t1630 259.26
R663 VDD.t2123 VDD.t2418 259.26
R664 VDD.t1299 VDD.t2123 259.26
R665 VDD.t2701 VDD.t1299 259.26
R666 VDD.t2552 VDD.t2701 259.26
R667 VDD.t990 VDD.t2552 259.26
R668 VDD.t2106 VDD.t990 259.26
R669 VDD.t3764 VDD.t2106 259.26
R670 VDD.t969 VDD.t3009 259.26
R671 VDD.t3009 VDD.t3945 259.26
R672 VDD.t3945 VDD.t2178 259.26
R673 VDD.t1999 VDD.t1822 259.26
R674 VDD.t1994 VDD.t1820 259.26
R675 VDD.t1996 VDD.t1818 259.26
R676 VDD.t1814 VDD.t1816 259.26
R677 VDD.t183 VDD.t179 259.26
R678 VDD.t607 VDD.t599 259.26
R679 VDD.t83 VDD.t1171 259.26
R680 VDD.t71 VDD.t69 259.26
R681 VDD.t63 VDD.t65 259.26
R682 VDD.t1326 VDD.t2880 259.26
R683 VDD.n1089 VDD.t4066 259.26
R684 VDD.t1243 VDD.n1089 259.26
R685 VDD.t1052 VDD.t1050 259.26
R686 VDD.t303 VDD.t309 259.26
R687 VDD.t311 VDD.t315 259.26
R688 VDD.n1957 VDD.t2142 259.26
R689 VDD.t2853 VDD.t494 259.26
R690 VDD.n915 VDD.t3684 259.26
R691 VDD.t3457 VDD.n915 259.26
R692 VDD.t2309 VDD.t878 259.26
R693 VDD.t3703 VDD.t2088 259.26
R694 VDD.t3982 VDD.t645 259.26
R695 VDD.t2003 VDD.t1920 259.26
R696 VDD.t1873 VDD.t1877 259.26
R697 VDD.t3501 VDD.t2428 259.26
R698 VDD.t1337 VDD.n238 259.26
R699 VDD.n238 VDD.t1054 259.26
R700 VDD.t4242 VDD.t4244 259.26
R701 VDD.t4246 VDD.t4248 259.26
R702 VDD.t1012 VDD.t1016 259.26
R703 VDD.t1004 VDD.t1006 259.26
R704 VDD.t1018 VDD.t1010 259.26
R705 VDD.t1008 VDD.t1014 259.26
R706 VDD.t2796 VDD.t2455 259.26
R707 VDD.t2837 VDD.t2796 259.26
R708 VDD.t2487 VDD.t2837 259.26
R709 VDD.t4236 VDD.t2487 259.26
R710 VDD.t2115 VDD.t4236 259.26
R711 VDD.t3301 VDD.t2115 259.26
R712 VDD.t3875 VDD.t3301 259.26
R713 VDD.t1441 VDD.t3875 259.26
R714 VDD.t3706 VDD.t3807 259.26
R715 VDD.t1559 VDD.t3706 259.26
R716 VDD.t1457 VDD.t1559 259.26
R717 VDD.t1515 VDD.t1457 259.26
R718 VDD.t1561 VDD.t1515 259.26
R719 VDD.t3396 VDD.t1561 259.26
R720 VDD.t3856 VDD.t3396 259.26
R721 VDD.t2597 VDD.t3856 259.26
R722 VDD.t2387 VDD.t2597 259.26
R723 VDD.t3889 VDD.t2387 259.26
R724 VDD.t3491 VDD.t3889 259.26
R725 VDD.t1147 VDD.t3491 259.26
R726 VDD.t4048 VDD.t1147 259.26
R727 VDD.t3210 VDD.t900 259.26
R728 VDD.t1188 VDD.t3210 259.26
R729 VDD.t951 VDD.t1188 259.26
R730 VDD.t3813 VDD.t951 259.26
R731 VDD.t1618 VDD.t3813 259.26
R732 VDD.t2305 VDD.t1618 259.26
R733 VDD.t2317 VDD.t2305 259.26
R734 VDD.t3927 VDD.t2317 259.26
R735 VDD.t3978 VDD.t3927 259.26
R736 VDD.t4160 VDD.t3978 259.26
R737 VDD.t3725 VDD.t4160 259.26
R738 VDD.t949 VDD.t3725 259.26
R739 VDD.t3565 VDD.t949 259.26
R740 VDD.t2155 VDD.t3565 259.26
R741 VDD.t2644 VDD.t2155 259.26
R742 VDD.t4015 VDD.t2644 259.26
R743 VDD.t2046 VDD.t2236 259.26
R744 VDD.t2067 VDD.t1401 259.26
R745 VDD.t3325 VDD.t2067 259.26
R746 VDD.t2378 VDD.t3325 259.26
R747 VDD.t2166 VDD.t2378 259.26
R748 VDD.t4264 VDD.t2166 259.26
R749 VDD.t1863 VDD.t4264 259.26
R750 VDD.t3271 VDD.t1863 259.26
R751 VDD.t2069 VDD.t3271 259.26
R752 VDD.t1521 VDD.t2069 259.26
R753 VDD.t1405 VDD.t1521 259.26
R754 VDD.t1169 VDD.t1405 259.26
R755 VDD.t4253 VDD.t1169 259.26
R756 VDD.t2772 VDD.t4253 259.26
R757 VDD.t2995 VDD.t2772 259.26
R758 VDD.t4003 VDD.t2995 259.26
R759 VDD.n2279 VDD.n2278 259.26
R760 VDD.t2017 VDD.t3148 259.26
R761 VDD.t2770 VDD.t2017 259.26
R762 VDD.t4278 VDD.t2770 259.26
R763 VDD.t2205 VDD.t4278 259.26
R764 VDD.t3997 VDD.t2205 259.26
R765 VDD.t1216 VDD.t3997 259.26
R766 VDD.t4255 VDD.t1216 259.26
R767 VDD.t2196 VDD.t4255 259.26
R768 VDD.t1763 VDD.t2585 259.26
R769 VDD.t4074 VDD.t1763 259.26
R770 VDD.t888 VDD.t882 259.26
R771 VDD.t884 VDD.t886 259.26
R772 VDD.t655 VDD.t629 259.26
R773 VDD.t623 VDD.t625 259.26
R774 VDD.t665 VDD.t653 259.26
R775 VDD.t627 VDD.t657 259.26
R776 VDD.t1513 VDD.t2745 258.065
R777 VDD.t2384 VDD.t2972 255.787
R778 VDD.t639 VDD.t1771 255.787
R779 VDD.t4061 VDD.t3858 255.787
R780 VDD.t895 VDD.t731 255.787
R781 VDD.t1160 VDD.t3460 253.472
R782 VDD.t846 VDD.t2647 253.472
R783 VDD.t3955 VDD.t3675 253.472
R784 VDD.t432 VDD.t769 251.157
R785 VDD.n1346 VDD.t2577 251.157
R786 VDD.t2847 VDD.t1278 251.087
R787 VDD.t434 VDD.t3958 250.299
R788 VDD.t835 VDD.t165 250
R789 VDD.t839 VDD.t163 250
R790 VDD.t833 VDD.t159 250
R791 VDD.t831 VDD.t161 250
R792 VDD.t287 VDD.t2751 250
R793 VDD.t1578 VDD.t3526 248.844
R794 VDD.t3931 VDD.t3933 247.685
R795 VDD.t725 VDD.t1508 247.685
R796 VDD.t3066 VDD.t3064 247.685
R797 VDD.t2960 VDD.t1848 244.214
R798 VDD.t4135 VDD.t3547 244.214
R799 VDD.t663 VDD.t3959 244.214
R800 VDD.t3618 VDD.t3622 243.728
R801 VDD.t1497 VDD.t3089 243.728
R802 VDD.t631 VDD.t775 243.728
R803 VDD.t860 VDD.t1894 243.148
R804 VDD.t2355 VDD.t3892 243.148
R805 VDD.t32 VDD.t37 243.148
R806 VDD.t617 VDD.t1084 243.148
R807 VDD.n401 VDD.t185 243.056
R808 VDD.t1960 VDD.t1209 243.056
R809 VDD.t1529 VDD.t2978 241.899
R810 VDD.t1512 VDD.t4300 241.899
R811 VDD.t2689 VDD.t3222 240.742
R812 VDD.t283 VDD.t289 240.742
R813 VDD.t1644 VDD.t2737 240.742
R814 VDD.t1896 VDD.t733 240.113
R815 VDD.t4230 VDD.t504 240.113
R816 VDD.t420 VDD.t426 239.897
R817 VDD.t3907 VDD.t2513 239.328
R818 VDD.t3570 VDD.t2097 238.427
R819 VDD.t1403 VDD.t1541 238.427
R820 VDD.t1266 VDD.t2240 238.389
R821 VDD.t30 VDD.t3394 237.978
R822 VDD.t721 VDD.t2074 237.269
R823 VDD.t1364 VDD.t1428 236.112
R824 VDD.t1366 VDD.t396 236.112
R825 VDD.t1112 VDD.t1611 236.112
R826 VDD.t3433 VDD.t1427 236.112
R827 VDD.t3604 VDD.t1111 236.112
R828 VDD.t1781 VDD.t4125 236.112
R829 VDD.t13 VDD.t693 236.112
R830 VDD.t4123 VDD.t1566 236.112
R831 VDD.t1565 VDD.t1407 236.112
R832 VDD.t779 VDD.t5 236.112
R833 VDD.t1594 VDD.t437 236.112
R834 VDD.t4013 VDD.t2986 236.112
R835 VDD.t3307 VDD.t4013 236.112
R836 VDD.t3033 VDD.t4262 236.112
R837 VDD.t17 VDD.t691 236.112
R838 VDD.t3216 VDD.t3281 236.112
R839 VDD.t1828 VDD.t4014 236.112
R840 VDD.t2470 VDD.t3217 236.112
R841 VDD.t3217 VDD.t948 236.112
R842 VDD.t3360 VDD.t2892 236.112
R843 VDD.t3710 VDD.t3361 236.112
R844 VDD.t358 VDD.t3358 236.112
R845 VDD.t3507 VDD.t531 236.112
R846 VDD.t944 VDD.t2742 236.112
R847 VDD.t2226 VDD.t1939 236.112
R848 VDD.t509 VDD.t2353 236.112
R849 VDD.t2052 VDD.t442 236.112
R850 VDD.t943 VDD.t3019 236.112
R851 VDD.t28 VDD.t2687 236.112
R852 VDD.t3819 VDD.t2406 236.112
R853 VDD.t3327 VDD.t3891 236.112
R854 VDD.t3023 VDD.t3388 236.112
R855 VDD.t3471 VDD.t3230 236.112
R856 VDD.t3479 VDD.t1808 236.112
R857 VDD.t3265 VDD.t1714 236.112
R858 VDD.t398 VDD.t1716 236.112
R859 VDD.t1075 VDD.t1090 236.112
R860 VDD.t3021 VDD.t3817 236.112
R861 VDD.t1527 VDD.t2814 236.112
R862 VDD.t819 VDD.t817 236.112
R863 VDD.t2813 VDD.t39 236.112
R864 VDD.t1079 VDD.t2813 236.112
R865 VDD.t35 VDD.t1079 236.112
R866 VDD.t3390 VDD.t35 236.112
R867 VDD.t4022 VDD.t475 236.112
R868 VDD.t3496 VDD.t2999 236.112
R869 VDD.t3072 VDD.t3496 236.112
R870 VDD.t1525 VDD.t3072 236.112
R871 VDD.t364 VDD.t3494 236.112
R872 VDD.t2906 VDD.t523 236.112
R873 VDD.t1966 VDD.t275 236.112
R874 VDD.t687 VDD.t699 236.112
R875 VDD.t4045 VDD.t1492 236.112
R876 VDD.t499 VDD.t2382 236.112
R877 VDD.t2268 VDD.t1035 236.112
R878 VDD.t823 VDD.t815 236.112
R879 VDD.t3785 VDD.t3954 236.112
R880 VDD.t2922 VDD.t3785 236.112
R881 VDD.t3489 VDD.t1095 236.112
R882 VDD.t1771 VDD.t4109 236.112
R883 VDD.t3858 VDD.t1066 236.112
R884 VDD.t3864 VDD.t3825 236.112
R885 VDD.t1056 VDD.t3860 236.112
R886 VDD.t651 VDD.t1056 236.112
R887 VDD.t1879 VDD.t3366 236.112
R888 VDD.t1203 VDD.t412 236.112
R889 VDD.t2948 VDD.t3583 236.112
R890 VDD.t2562 VDD.t2311 236.112
R891 VDD.t1092 VDD.t787 236.112
R892 VDD.t3815 VDD.t963 236.112
R893 VDD.t1773 VDD.t3815 236.112
R894 VDD.t1279 VDD.t2080 236.112
R895 VDD.t3582 VDD.t4007 236.112
R896 VDD.t9 VDD.t895 236.112
R897 VDD.t3466 VDD.t729 236.112
R898 VDD.t1519 VDD.t3749 236.112
R899 VDD.t0 VDD.t2191 236.112
R900 VDD.t494 VDD.t3887 236.112
R901 VDD.t2543 VDD.t1838 236.112
R902 VDD.t2412 VDD.t3722 236.112
R903 VDD.t3722 VDD.t897 236.112
R904 VDD.t2620 VDD.t1506 236.112
R905 VDD.t1672 VDD.t2083 236.112
R906 VDD.t3848 VDD.t2141 236.112
R907 VDD.t3920 VDD.t1962 236.112
R908 VDD.t3597 VDD.t3150 236.112
R909 VDD.t3991 VDD.t1413 236.112
R910 VDD.t1453 VDD.t2035 236.112
R911 VDD.t1648 VDD.t2285 236.112
R912 VDD.t1638 VDD.t1646 236.112
R913 VDD.t1642 VDD.t1650 236.112
R914 VDD.t1640 VDD.t1636 236.112
R915 VDD.t761 VDD.t2734 236.112
R916 VDD.t771 VDD.t715 236.112
R917 VDD.t2257 VDD.t648 236.112
R918 VDD.t3273 VDD.t3490 236.112
R919 VDD.t2238 VDD.t4107 236.112
R920 VDD.t488 VDD.t1908 236.112
R921 VDD.t1454 VDD.t2827 236.112
R922 VDD.t2747 VDD.t1382 235.963
R923 VDD.t1268 VDD.t2763 234.954
R924 VDD.t1146 VDD.t1998 234.954
R925 VDD.t2786 VDD.t2706 234.625
R926 VDD.t1062 VDD.n432 233.797
R927 VDD.t1038 VDD.t2054 233.612
R928 VDD.t1386 VDD.t1380 233.061
R929 VDD.t1973 VDD.t2930 232.639
R930 VDD.t2862 VDD.t3606 232.639
R931 VDD.t2924 VDD.n2023 232.639
R932 VDD.t4122 VDD.t634 232.639
R933 VDD.t3363 VDD.t1670 232.274
R934 VDD.t2140 VDD.t3743 232.274
R935 VDD.t3051 VDD.t2983 231.685
R936 VDD.t335 VDD.t4092 231.482
R937 VDD.t920 VDD.t2950 231.482
R938 VDD.t910 VDD.t85 231.482
R939 VDD.t2176 VDD.t307 231.482
R940 VDD.t1533 VDD.t1918 231.482
R941 VDD.t1830 VDD.t3493 230.585
R942 VDD.t4070 VDD.t3951 230.585
R943 VDD.t2976 VDD.t3447 230.325
R944 VDD.t2222 VDD.t3083 230.325
R945 VDD.t1836 VDD.t485 230.325
R946 VDD.t277 VDD.t1276 229.77
R947 VDD.t422 VDD.t1000 228.01
R948 VDD.t3415 VDD.t2497 228.01
R949 VDD.t1702 VDD.t2920 228.01
R950 VDD.t4114 VDD.t3256 228.01
R951 VDD.t1892 VDD.t1859 228.01
R952 VDD.t2512 VDD.t3901 226.852
R953 VDD.t1430 VDD.t1360 226.852
R954 VDD.t3228 VDD.t4086 226.852
R955 VDD.t3039 VDD.t2019 226.852
R956 VDD.t829 VDD.t169 226.852
R957 VDD.t827 VDD.t167 226.852
R958 VDD.t837 VDD.t157 226.852
R959 VDD.t841 VDD.t187 226.852
R960 VDD.t1806 VDD.t141 226.852
R961 VDD.t1968 VDD.t151 226.852
R962 VDD.t916 VDD.t2268 226.852
R963 VDD.t1033 VDD.t2532 226.852
R964 VDD.t492 VDD.t441 226.852
R965 VDD.t726 VDD.t1365 226.394
R966 VDD.t2908 VDD.t3661 225.695
R967 VDD.t778 VDD.t784 225.695
R968 VDD.t501 VDD.t2376 225.695
R969 VDD.t3127 VDD.t1729 225.695
R970 VDD.t536 VDD.t488 225.695
R971 VDD.t205 VDD.t2544 225.695
R972 VDD.t362 VDD.n517 224.537
R973 VDD.t3911 VDD.t2764 224.537
R974 VDD.n1950 VDD.t2618 224.537
R975 VDD.t533 VDD.t3669 223.716
R976 VDD.t465 VDD.t2989 223.716
R977 VDD.t424 VDD.t3646 223.381
R978 VDD.t3750 VDD.t3047 223.381
R979 VDD.t2866 VDD.t539 223.381
R980 VDD.t2184 VDD.t2332 222.222
R981 VDD.t1263 VDD.t852 222.222
R982 VDD.t1963 VDD.t2948 222.222
R983 VDD.t4044 VDD.t1257 221.065
R984 VDD.t1826 VDD.t739 219.907
R985 VDD.t704 VDD.t3283 219.907
R986 VDD.t11 VDD.t1660 219.907
R987 VDD.t3542 VDD.n1604 218.75
R988 VDD.t3017 VDD.n1597 218.75
R989 VDD.t1859 VDD.n441 218.75
R990 VDD.t2952 VDD.n1788 218.75
R991 VDD.t992 VDD.n1957 218.75
R992 VDD.t1571 VDD.n269 218.75
R993 VDD.t946 VDD.t3214 217.594
R994 VDD.t3488 VDD.t3331 217.594
R995 VDD.t67 VDD.t2136 217.594
R996 VDD.t301 VDD.t1120 217.594
R997 VDD.t2001 VDD.t3850 217.594
R998 VDD.t2426 VDD.t507 217.594
R999 VDD.n1393 VDD.t2470 215.279
R1000 VDD.t1556 VDD.t1550 215.279
R1001 VDD.t1965 VDD.t697 215.054
R1002 VDD.t765 VDD.t3138 214.444
R1003 VDD.t2687 VDD.t537 214.444
R1004 VDD.t3919 VDD.n262 214.12
R1005 VDD.t3393 VDD.t603 212.964
R1006 VDD.t2819 VDD.t1552 212.964
R1007 VDD.t3679 VDD.t19 212.964
R1008 VDD.t643 VDD.t1337 212.964
R1009 VDD.t777 VDD.t3200 212.964
R1010 VDD.t3700 VDD.t3386 212.964
R1011 VDD.t1173 VDD.t1493 212.143
R1012 VDD.t313 VDD.t1093 212.143
R1013 VDD.t1875 VDD.t3791 212.143
R1014 VDD.t4009 VDD.t723 211.806
R1015 VDD.t3028 VDD.t2 210.649
R1016 VDD.t279 VDD.t3339 209.913
R1017 VDD.t3413 VDD.t1376 209.492
R1018 VDD.t1951 VDD.t4165 209.492
R1019 VDD.t2946 VDD.t3471 209.492
R1020 VDD.t2088 VDD.t4299 209.492
R1021 VDD.t1834 VDD.t3355 209.492
R1022 VDD.t2480 VDD.t2078 209.081
R1023 VDD.t3909 VDD.t708 208.333
R1024 VDD.t1895 VDD.t3659 208.333
R1025 VDD.t1027 VDD.t2518 208.333
R1026 VDD.t1166 VDD.t4094 208.333
R1027 VDD.t2882 VDD.t821 208.333
R1028 VDD.t147 VDD.t177 208.333
R1029 VDD.t145 VDD.t171 208.333
R1030 VDD.t3630 VDD.t1295 208.333
R1031 VDD.t3355 VDD.t2412 208.333
R1032 VDD.t3766 VDD.t783 207.177
R1033 VDD.t2428 VDD.t2257 207.177
R1034 VDD.t1959 VDD.t2258 206.691
R1035 VDD.t3140 VDD.t1429 206.019
R1036 VDD.t1869 VDD.t2914 204.862
R1037 VDD.t1230 VDD.t3254 204.862
R1038 VDD.t880 VDD.t3066 204.862
R1039 VDD.t902 VDD.t3895 203.704
R1040 VDD.t3993 VDD.t850 203.704
R1041 VDD.t295 VDD.t4261 203.704
R1042 VDD.t299 VDD.t1286 203.704
R1043 VDD.t410 VDD.t1463 203.704
R1044 VDD.t439 VDD.t3474 203.704
R1045 VDD.t3402 VDD.t767 202.547
R1046 VDD.t4024 VDD.t3604 202.547
R1047 VDD.t2198 VDD.t3540 202.547
R1048 VDD.t711 VDD.t749 202.547
R1049 VDD.t1861 VDD.t3498 202.547
R1050 VDD.t34 VDD.t802 202.308
R1051 VDD.t1128 VDD.n577 201.389
R1052 VDD.t195 VDD.n600 201.389
R1053 VDD.t3797 VDD.t3293 201.389
R1054 VDD.n1597 VDD.t7 201.389
R1055 VDD.t1155 VDD.t2180 201.389
R1056 VDD.n1788 VDD.t1891 201.389
R1057 VDD.t599 VDD.n1775 201.389
R1058 VDD.t788 VDD.n1950 201.389
R1059 VDD.t1838 VDD.t3692 201.389
R1060 VDD.t4300 VDD.t3982 201.389
R1061 VDD.t1211 VDD.t3920 201.389
R1062 VDD.t1140 VDD.t3487 201.389
R1063 VDD.t1726 VDD.t4078 201.389
R1064 VDD.t1791 VDD.t2033 201.389
R1065 VDD.t3125 VDD.n2104 201.389
R1066 VDD.t3716 VDD.n2174 201.389
R1067 VDD.t4248 VDD.t2400 201.389
R1068 VDD.t1016 VDD.t4268 201.389
R1069 VDD.t1006 VDD.t1933 201.389
R1070 VDD.t1010 VDD.t2884 201.389
R1071 VDD.t1014 VDD.t4051 201.389
R1072 VDD.t882 VDD.t4074 201.389
R1073 VDD.t886 VDD.t1205 201.389
R1074 VDD.t629 VDD.t3226 201.389
R1075 VDD.t625 VDD.t2938 201.389
R1076 VDD.t653 VDD.t1851 201.389
R1077 VDD.t657 VDD.t4099 201.389
R1078 VDD.t1374 VDD.t1720 200.718
R1079 VDD.t1958 VDD.t1956 200.718
R1080 VDD.t1193 VDD.t1192 200.718
R1081 VDD.t3481 VDD.t3482 200.238
R1082 VDD.t2616 VDD.t4205 199.075
R1083 VDD.t3560 VDD.t3909 198.254
R1084 VDD.t659 VDD.t1807 197.917
R1085 VDD.t4220 VDD.t2108 196.76
R1086 VDD.t3189 VDD.t2389 196.76
R1087 VDD.t1767 VDD.t20 195.602
R1088 VDD.t2970 VDD.t3104 194.744
R1089 VDD.t428 VDD.t754 194.445
R1090 VDD.t4251 VDD.t4250 194.445
R1091 VDD.t3322 VDD.t3324 194.445
R1092 VDD.t2649 VDD.t2650 194.445
R1093 VDD.t1848 VDD.t1850 194.445
R1094 VDD.t4036 VDD.t4035 194.445
R1095 VDD.t3780 VDD.t3782 194.445
R1096 VDD.t3116 VDD.t3114 194.445
R1097 VDD.t4224 VDD.t4222 194.445
R1098 VDD.t1711 VDD.t1709 194.445
R1099 VDD.t3547 VDD.t3546 194.445
R1100 VDD.t2131 VDD.t2133 194.445
R1101 VDD.t1950 VDD.t1951 194.445
R1102 VDD.t1349 VDD.t1347 194.445
R1103 VDD.t2763 VDD.t2761 194.445
R1104 VDD.t2748 VDD.t2750 194.445
R1105 VDD.t1808 VDD.t1449 194.445
R1106 VDD.t1399 VDD.t1398 194.445
R1107 VDD.t638 VDD.t3299 194.445
R1108 VDD.t2568 VDD.t2566 194.445
R1109 VDD.t1144 VDD.t1146 194.445
R1110 VDD.t2165 VDD.t2163 194.445
R1111 VDD.t477 VDD.t1173 194.445
R1112 VDD.t2880 VDD.t2879 194.445
R1113 VDD.t1113 VDD.t1114 194.445
R1114 VDD.t1284 VDD.t297 194.445
R1115 VDD.t3519 VDD.t3517 194.445
R1116 VDD.t2212 VDD.t2211 194.445
R1117 VDD.t4209 VDD.t3864 194.445
R1118 VDD.t517 VDD.t313 194.445
R1119 VDD.t3177 VDD.t3175 194.445
R1120 VDD.t3184 VDD.t3186 194.445
R1121 VDD.t4299 VDD.t4297 194.445
R1122 VDD.t497 VDD.t1875 194.445
R1123 VDD.t1184 VDD.t1183 194.445
R1124 VDD.t1881 VDD.t1883 194.445
R1125 VDD.t3357 VDD.t2199 193.548
R1126 VDD.t1074 VDD.t1925 193.287
R1127 VDD.t605 VDD.t7 193.287
R1128 VDD.t2918 VDD.t2689 193.287
R1129 VDD.n473 VDD.t3925 193.287
R1130 VDD.t1199 VDD.t1994 193.287
R1131 VDD.t289 VDD.t3755 193.287
R1132 VDD.t717 VDD.t2784 192.131
R1133 VDD.t3285 VDD.t3218 192.131
R1134 VDD.t238 VDD.n334 192.131
R1135 VDD.t921 VDD.t3073 191.756
R1136 VDD.t374 VDD.t372 191.388
R1137 VDD.t378 VDD.t374 191.388
R1138 VDD.t380 VDD.t378 191.388
R1139 VDD.t384 VDD.t380 191.388
R1140 VDD.t368 VDD.t384 191.388
R1141 VDD.t382 VDD.t368 191.388
R1142 VDD.t366 VDD.t382 191.388
R1143 VDD.t370 VDD.t366 191.388
R1144 VDD.t376 VDD.t370 191.388
R1145 VDD.t339 VDD.t341 191.388
R1146 VDD.t341 VDD.t337 191.388
R1147 VDD.t337 VDD.t343 191.388
R1148 VDD.t343 VDD.t345 191.388
R1149 VDD.t345 VDD.t325 191.388
R1150 VDD.t325 VDD.t327 191.388
R1151 VDD.t327 VDD.t333 191.388
R1152 VDD.t333 VDD.t329 191.388
R1153 VDD.t329 VDD.t331 191.388
R1154 VDD.t206 VDD.t214 191.388
R1155 VDD.t212 VDD.t206 191.388
R1156 VDD.t209 VDD.t212 191.388
R1157 VDD.t215 VDD.t209 191.388
R1158 VDD.t211 VDD.t215 191.388
R1159 VDD.t208 VDD.t211 191.388
R1160 VDD.t210 VDD.t208 191.388
R1161 VDD.t207 VDD.t210 191.388
R1162 VDD.t213 VDD.t207 191.388
R1163 VDD.t232 VDD.t220 191.388
R1164 VDD.t224 VDD.t232 191.388
R1165 VDD.t218 VDD.t224 191.388
R1166 VDD.t230 VDD.t218 191.388
R1167 VDD.t216 VDD.t230 191.388
R1168 VDD.t228 VDD.t216 191.388
R1169 VDD.t222 VDD.t228 191.388
R1170 VDD.t234 VDD.t222 191.388
R1171 VDD.t226 VDD.t234 191.388
R1172 VDD.t1903 VDD.t1847 191.388
R1173 VDD.t1845 VDD.t1903 191.388
R1174 VDD.t1842 VDD.t1845 191.388
R1175 VDD.t1902 VDD.t1842 191.388
R1176 VDD.t1844 VDD.t1902 191.388
R1177 VDD.t1905 VDD.t1844 191.388
R1178 VDD.t1843 VDD.t1905 191.388
R1179 VDD.t1904 VDD.t1843 191.388
R1180 VDD.t1846 VDD.t1904 191.388
R1181 VDD.t593 VDD.t581 191.388
R1182 VDD.t585 VDD.t593 191.388
R1183 VDD.t579 VDD.t585 191.388
R1184 VDD.t591 VDD.t579 191.388
R1185 VDD.t577 VDD.t591 191.388
R1186 VDD.t589 VDD.t577 191.388
R1187 VDD.t583 VDD.t589 191.388
R1188 VDD.t595 VDD.t583 191.388
R1189 VDD.t587 VDD.t595 191.388
R1190 VDD.t2694 VDD.t2699 191.388
R1191 VDD.t2697 VDD.t2694 191.388
R1192 VDD.t2700 VDD.t2697 191.388
R1193 VDD.t2693 VDD.t2700 191.388
R1194 VDD.t2696 VDD.t2693 191.388
R1195 VDD.t2691 VDD.t2696 191.388
R1196 VDD.t2695 VDD.t2691 191.388
R1197 VDD.t2698 VDD.t2695 191.388
R1198 VDD.t2692 VDD.t2698 191.388
R1199 VDD.t567 VDD.t555 191.388
R1200 VDD.t551 VDD.t567 191.388
R1201 VDD.t559 VDD.t551 191.388
R1202 VDD.t565 VDD.t559 191.388
R1203 VDD.t553 VDD.t565 191.388
R1204 VDD.t563 VDD.t553 191.388
R1205 VDD.t569 VDD.t563 191.388
R1206 VDD.t557 VDD.t569 191.388
R1207 VDD.t561 VDD.t557 191.388
R1208 VDD.t107 VDD.t112 191.388
R1209 VDD.t110 VDD.t107 191.388
R1210 VDD.t113 VDD.t110 191.388
R1211 VDD.t116 VDD.t113 191.388
R1212 VDD.t109 VDD.t116 191.388
R1213 VDD.t114 VDD.t109 191.388
R1214 VDD.t108 VDD.t114 191.388
R1215 VDD.t111 VDD.t108 191.388
R1216 VDD.t115 VDD.t111 191.388
R1217 VDD.t679 VDD.t667 191.388
R1218 VDD.t683 VDD.t679 191.388
R1219 VDD.t671 VDD.t683 191.388
R1220 VDD.t677 VDD.t671 191.388
R1221 VDD.t685 VDD.t677 191.388
R1222 VDD.t675 VDD.t685 191.388
R1223 VDD.t681 VDD.t675 191.388
R1224 VDD.t669 VDD.t681 191.388
R1225 VDD.t673 VDD.t669 191.388
R1226 VDD.t547 VDD.t542 191.388
R1227 VDD.t550 VDD.t547 191.388
R1228 VDD.t543 VDD.t550 191.388
R1229 VDD.t546 VDD.t543 191.388
R1230 VDD.t549 VDD.t546 191.388
R1231 VDD.t544 VDD.t549 191.388
R1232 VDD.t548 VDD.t544 191.388
R1233 VDD.t541 VDD.t548 191.388
R1234 VDD.t545 VDD.t541 191.388
R1235 VDD.t255 VDD.t263 191.388
R1236 VDD.t259 VDD.t255 191.388
R1237 VDD.t267 VDD.t259 191.388
R1238 VDD.t253 VDD.t267 191.388
R1239 VDD.t261 VDD.t253 191.388
R1240 VDD.t271 VDD.t261 191.388
R1241 VDD.t257 VDD.t271 191.388
R1242 VDD.t265 VDD.t257 191.388
R1243 VDD.t269 VDD.t265 191.388
R1244 VDD.t133 VDD.t131 191.388
R1245 VDD.t129 VDD.t133 191.388
R1246 VDD.t136 VDD.t129 191.388
R1247 VDD.t132 VDD.t136 191.388
R1248 VDD.t128 VDD.t132 191.388
R1249 VDD.t135 VDD.t128 191.388
R1250 VDD.t127 VDD.t135 191.388
R1251 VDD.t134 VDD.t127 191.388
R1252 VDD.t130 VDD.t134 191.388
R1253 VDD.t1749 VDD.t1757 191.388
R1254 VDD.t1741 VDD.t1749 191.388
R1255 VDD.t1755 VDD.t1741 191.388
R1256 VDD.t1747 VDD.t1755 191.388
R1257 VDD.t1753 VDD.t1747 191.388
R1258 VDD.t1745 VDD.t1753 191.388
R1259 VDD.t1759 VDD.t1745 191.388
R1260 VDD.t1751 VDD.t1759 191.388
R1261 VDD.t1743 VDD.t1751 191.388
R1262 VDD.t79 VDD.t77 191.388
R1263 VDD.t75 VDD.t79 191.388
R1264 VDD.t82 VDD.t75 191.388
R1265 VDD.t78 VDD.t82 191.388
R1266 VDD.t74 VDD.t78 191.388
R1267 VDD.t81 VDD.t74 191.388
R1268 VDD.t73 VDD.t81 191.388
R1269 VDD.t80 VDD.t73 191.388
R1270 VDD.t76 VDD.t80 191.388
R1271 VDD.t1303 VDD.t1311 191.388
R1272 VDD.t1315 VDD.t1303 191.388
R1273 VDD.t1309 VDD.t1315 191.388
R1274 VDD.t1301 VDD.t1309 191.388
R1275 VDD.t1307 VDD.t1301 191.388
R1276 VDD.t1319 VDD.t1307 191.388
R1277 VDD.t1313 VDD.t1319 191.388
R1278 VDD.t1305 VDD.t1313 191.388
R1279 VDD.t1317 VDD.t1305 191.388
R1280 VDD.t404 VDD.t402 191.388
R1281 VDD.t400 VDD.t404 191.388
R1282 VDD.t407 VDD.t400 191.388
R1283 VDD.t403 VDD.t407 191.388
R1284 VDD.t409 VDD.t403 191.388
R1285 VDD.t406 VDD.t409 191.388
R1286 VDD.t408 VDD.t406 191.388
R1287 VDD.t405 VDD.t408 191.388
R1288 VDD.t401 VDD.t405 191.388
R1289 VDD.t89 VDD.t97 191.388
R1290 VDD.t101 VDD.t89 191.388
R1291 VDD.t95 VDD.t101 191.388
R1292 VDD.t87 VDD.t95 191.388
R1293 VDD.t93 VDD.t87 191.388
R1294 VDD.t105 VDD.t93 191.388
R1295 VDD.t99 VDD.t105 191.388
R1296 VDD.t91 VDD.t99 191.388
R1297 VDD.t103 VDD.t91 191.388
R1298 VDD.t1261 VDD.t4216 190.972
R1299 VDD.t3224 VDD.t609 189.815
R1300 VDD.t4127 VDD.t819 189.815
R1301 VDD.t4195 VDD.t3123 189.815
R1302 VDD.t1824 VDD.t55 187.5
R1303 VDD.t2581 VDD.t2501 187.5
R1304 VDD.n1393 VDD.t946 187.5
R1305 VDD.t1029 VDD.n494 187.5
R1306 VDD.t1820 VDD.t1451 187.5
R1307 VDD.t1818 VDD.t2573 187.5
R1308 VDD.t3921 VDD.t430 186.381
R1309 VDD.t20 VDD.t4251 186.344
R1310 VDD.t1036 VDD.t183 186.344
R1311 VDD.t3186 VDD.t2309 186.344
R1312 VDD.t449 VDD.t2293 185.185
R1313 VDD.t1372 VDD.t4018 185.185
R1314 VDD.t1563 VDD.t3663 185.185
R1315 VDD.t3260 VDD.t615 185.185
R1316 VDD.t2109 VDD.t4147 185.185
R1317 VDD.t2108 VDD.t4148 185.185
R1318 VDD.t2508 VDD.t3189 185.185
R1319 VDD.t2507 VDD.t3190 185.185
R1320 VDD.t4088 VDD.t2326 185.185
R1321 VDD.t153 VDD.t175 185.185
R1322 VDD.t149 VDD.t173 185.185
R1323 VDD.t2588 VDD.t486 185.185
R1324 VDD.t733 VDD.t61 184.744
R1325 VDD.t2328 VDD.t944 184.029
R1326 VDD.t739 VDD.t1712 182.87
R1327 VDD.t1181 VDD.t704 182.87
R1328 VDD.t1237 VDD.t317 182.87
R1329 VDD.t473 VDD.t533 182.87
R1330 VDD.t2144 VDD.t2841 182.87
R1331 VDD.t2040 VDD.t2654 182.87
R1332 VDD.t483 VDD.t465 182.87
R1333 VDD.t1114 VDD.t4120 181.714
R1334 VDD.t3735 VDD.t2964 181.601
R1335 VDD.t37 VDD.t4026 181.168
R1336 VDD.t763 VDD.t1372 180.556
R1337 VDD.t3624 VDD.t1153 180.556
R1338 VDD.t2180 VDD.t3844 180.556
R1339 VDD.t2121 VDD.t143 180.556
R1340 VDD.t1220 VDD.t3096 180.556
R1341 VDD.t3475 VDD.t1963 180.556
R1342 VDD.t441 VDD.t4030 179.734
R1343 VDD.t4129 VDD.t2104 179.399
R1344 VDD.t3264 VDD.t1064 179.399
R1345 VDD.t3106 VDD.t3600 179.399
R1346 VDD.n420 VDD.t3553 179.212
R1347 VDD.t815 VDD.t758 178.242
R1348 VDD.t731 VDD.t4152 178.242
R1349 VDD.t22 VDD.t3505 178.018
R1350 VDD.n373 VDD.t440 177.226
R1351 VDD.t2225 VDD.t2671 176.822
R1352 VDD.t945 VDD.t2223 176.822
R1353 VDD.t2814 VDD.n420 176.226
R1354 VDD.t3437 VDD.t3957 175.927
R1355 VDD.t12 VDD.t3297 175.927
R1356 VDD.t2019 VDD.t2952 175.927
R1357 VDD.t3175 VDD.t2057 175.927
R1358 VDD.t2497 VDD.t1573 174.769
R1359 VDD.t861 VDD.t3657 174.769
R1360 VDD.t2015 VDD.t1892 174.769
R1361 VDD.t463 VDD.t1325 174.769
R1362 VDD.t1883 VDD.t3273 174.769
R1363 VDD.t1554 VDD.t727 173.612
R1364 VDD.t3954 VDD.t1267 173.612
R1365 VDD.t3569 VDD.t1735 173.612
R1366 VDD.t1948 VDD.t1543 173.612
R1367 VDD.t2191 VDD.t644 173.612
R1368 VDD.t2859 VDD.t2313 173.612
R1369 VDD.t1837 VDD.t2564 173.612
R1370 VDD.t3338 VDD.t3620 173.238
R1371 VDD.t4165 VDD.t3871 172.454
R1372 VDD.t506 VDD.t3192 172.454
R1373 VDD.t4297 VDD.t1834 172.454
R1374 VDD.t811 VDD.t1077 171.633
R1375 VDD.t1486 VDD.t191 171.297
R1376 VDD.t2768 VDD.t1656 171.297
R1377 VDD.t1407 VDD.t428 171.297
R1378 VDD.t1362 VDD.t2222 171.297
R1379 VDD.t1939 VDD.t3030 171.297
R1380 VDD.t2356 VDD.t1282 171.297
R1381 VDD.t1035 VDD.t1220 171.297
R1382 VDD.t1871 VDD.t790 171.297
R1383 VDD.t1470 VDD.t22 170.849
R1384 VDD.t2073 VDD.t1364 170.139
R1385 VDD.t796 VDD.t2408 170.139
R1386 VDD.t2930 VDD.t3542 170.139
R1387 VDD.t137 VDD.t1603 170.139
R1388 VDD.n2023 VDD.t3692 170.139
R1389 VDD.n303 VDD.t1505 168.982
R1390 VDD.t2461 VDD.t1356 168.982
R1391 VDD.t1729 VDD.n255 168.982
R1392 VDD.t2282 VDD.t718 168.982
R1393 VDD.t15 VDD.t771 167.825
R1394 VDD.t3553 VDD.t3735 167.264
R1395 VDD.t1597 VDD.t392 166.667
R1396 VDD.t1467 VDD.t1776 166.667
R1397 VDD.t864 VDD.t318 166.667
R1398 VDD.t2904 VDD.t3733 166.667
R1399 VDD.t65 VDD.t2626 166.667
R1400 VDD.t2740 VDD.t3952 166.667
R1401 VDD.t4284 VDD.t646 166.667
R1402 VDD.t2854 VDD.t2059 166.667
R1403 VDD.t3862 VDD.t601 165.51
R1404 VDD.t1068 VDD.t809 165.51
R1405 VDD.t3503 VDD.t3588 165.51
R1406 VDD.t3493 VDD.t921 163.68
R1407 VDD.t3951 VDD.t1931 163.68
R1408 VDD.t2535 VDD.t711 163.195
R1409 VDD.t3094 VDD.t181 163.195
R1410 VDD.t430 VDD.t1568 162.486
R1411 VDD.n348 VDD.t1795 162.099
R1412 VDD.t1378 VDD.t1783 162.037
R1413 VDD.t3361 VDD.t2788 162.037
R1414 VDD.t3222 VDD.t3840 162.037
R1415 VDD.t1867 VDD.t2924 162.037
R1416 VDD.n2115 VDD.n2114 161.236
R1417 VDD.t2723 VDD.t1527 160.881
R1418 VDD.t1168 VDD.t706 160.881
R1419 VDD.t2978 VDD.t2524 160.881
R1420 VDD.t24 VDD.t1529 160.881
R1421 VDD.t1048 VDD.t1531 160.881
R1422 VDD.t3138 VDD.t1352 159.722
R1423 VDD.t1209 VDD.t2466 159.722
R1424 VDD.t1795 VDD.t238 159.346
R1425 VDD.t285 VDD.t1255 157.407
R1426 VDD.t2532 VDD.n373 156.552
R1427 VDD.t1573 VDD.n610 156.25
R1428 VDD.t1066 VDD.t639 156.25
R1429 VDD.t3620 VDD.t2705 155.498
R1430 VDD.t649 VDD.t4061 155.094
R1431 VDD.t3985 VDD.t413 155.094
R1432 VDD.t3104 VDD.t1715 154.123
R1433 VDD.t735 VDD.t3433 153.935
R1434 VDD.t2133 VDD.t2410 153.935
R1435 VDD.t2080 VDD.t4009 153.935
R1436 VDD.t2223 VDD.t3216 153.733
R1437 VDD.t356 VDD.t2717 152.779
R1438 VDD.t1943 VDD.t193 152.779
R1439 VDD.t2974 VDD.t1654 152.779
R1440 VDD.t573 VDD.t3866 152.779
R1441 VDD.t117 VDD.t125 152.779
R1442 VDD.t121 VDD.t621 152.779
R1443 VDD.t319 VDD.t2608 152.779
R1444 VDD.t354 VDD.t2634 152.779
R1445 VDD.t347 VDD.t2614 152.779
R1446 VDD.t390 VDD.t2612 152.779
R1447 VDD.t1891 VDD.t1222 152.779
R1448 VDD.t275 VDD.t607 152.779
R1449 VDD.t3076 VDD.t2432 152.779
R1450 VDD.t1700 VDD.t744 151.62
R1451 VDD.t445 VDD.t4115 151.62
R1452 VDD.t1352 VDD.t2936 150.464
R1453 VDD.t2624 VDD.t4258 150.464
R1454 VDD.t3606 VDD.t1396 149.306
R1455 VDD.t1954 VDD.t1274 149.306
R1456 VDD.t1784 VDD.t1374 148.149
R1457 VDD.t352 VDD.t123 148.149
R1458 VDD.t2434 VDD.t2426 148.149
R1459 VDD.t800 VDD.t34 147.796
R1460 VDD.t3648 VDD.t1128 146.992
R1461 VDD.n1272 VDD.t1459 145.833
R1462 VDD.t1044 VDD.t4145 145.833
R1463 VDD.t2528 VDD.t4173 145.833
R1464 VDD.t2877 VDD.t1341 145.833
R1465 VDD.t1956 VDD.t3357 145.76
R1466 VDD.t2199 VDD.t3362 145.504
R1467 VDD.t3667 VDD.t721 144.677
R1468 VDD.t3801 VDD.t2186 144.677
R1469 VDD.t2731 VDD.t2170 144.677
R1470 VDD.t2311 VDD.t788 144.677
R1471 VDD.t3879 VDD.t3059 143.519
R1472 VDD.t1586 VDD.t862 143.519
R1473 VDD.t3259 VDD.t3220 143.519
R1474 VDD.t4145 VDD.t1046 143.519
R1475 VDD.t3024 VDD.t613 143.519
R1476 VDD.t4133 VDD.t1070 143.519
R1477 VDD.t807 VDD.t1042 143.519
R1478 VDD.t813 VDD.t26 143.519
R1479 VDD.t597 VDD.t1086 143.519
R1480 VDD.t1088 VDD.t1060 143.519
R1481 VDD.t2050 VDD.t1058 143.519
R1482 VDD.t3551 VDD.t825 143.519
R1483 VDD.t39 VDD.t3698 143.519
R1484 VDD.t4065 VDD.t1525 143.519
R1485 VDD.t416 VDD.t1490 143.519
R1486 VDD.t305 VDD.t3364 143.519
R1487 VDD.t2097 VDD.t3595 143.519
R1488 VDD.t2436 VDD.t1403 143.519
R1489 VDD.t1 VDD.t2587 143.519
R1490 VDD.t2005 VDD.t2138 143.519
R1491 VDD.t1624 VDD.t3612 143.519
R1492 VDD.t1855 VDD.t3446 142.362
R1493 VDD.t929 VDD.t2131 142.362
R1494 VDD.t1880 VDD.t1664 142.362
R1495 VDD.t3849 VDD.t3741 142.362
R1496 VDD.t4111 VDD.t2099 141.204
R1497 VDD.t3661 VDD.t1896 140.047
R1498 VDD.t1728 VDD.t2480 139.786
R1499 VDD.t1477 VDD.t687 139.5
R1500 VDD.t2258 VDD.t3919 139.036
R1501 VDD.t1384 VDD.t2746 138.889
R1502 VDD.t3444 VDD.t2541 138.889
R1503 VDD.t693 VDD.t195 137.732
R1504 VDD.t2161 VDD.t2960 137.732
R1505 VDD.t2577 VDD.t4135 137.732
R1506 VDD.t3925 VDD.t3720 137.732
R1507 VDD.t1870 VDD.t1062 137.732
R1508 VDD.t3757 VDD.t3823 137.732
R1509 VDD.t3817 VDD.t3731 137.732
R1510 VDD.t3212 VDD.t2076 137.732
R1511 VDD.t723 VDD.n1949 136.575
R1512 VDD.t1505 VDD.t323 136.575
R1513 VDD.t3511 VDD.t3017 135.417
R1514 VDD.t3758 VDD.t1334 135.417
R1515 VDD.t1118 VDD.t1052 135.417
R1516 VDD.t1287 VDD.t992 135.417
R1517 VDD.t3705 VDD.t877 135.417
R1518 VDD.t897 VDD.t636 135.417
R1519 VDD.t1601 VDD.t1565 134.26
R1520 VDD.t1109 VDD.t573 134.26
R1521 VDD.t3807 VDD.n650 133.941
R1522 VDD.t697 VDD.t1477 133.811
R1523 VDD.t744 VDD.t735 133.102
R1524 VDD.t1050 VDD.t1871 131.945
R1525 VDD.t2685 VDD.t3650 131.945
R1526 VDD.t4115 VDD.t823 130.787
R1527 VDD.t2397 VDD.t906 130.095
R1528 VDD.n1508 VDD.n560 129.631
R1529 VDD.t2715 VDD.t2514 129.631
R1530 VDD.t2514 VDD.t2713 129.631
R1531 VDD.t49 VDD.t251 129.631
R1532 VDD.t251 VDD.t51 129.631
R1533 VDD.t51 VDD.t273 129.631
R1534 VDD.t273 VDD.t59 129.631
R1535 VDD.t59 VDD.t245 129.631
R1536 VDD.t245 VDD.t47 129.631
R1537 VDD.t47 VDD.t249 129.631
R1538 VDD.t249 VDD.t870 129.631
R1539 VDD.t870 VDD.t241 129.631
R1540 VDD.t241 VDD.t866 129.631
R1541 VDD.t866 VDD.t243 129.631
R1542 VDD.t243 VDD.t872 129.631
R1543 VDD.t872 VDD.t247 129.631
R1544 VDD.t247 VDD.t868 129.631
R1545 VDD.t868 VDD.t239 129.631
R1546 VDD.t197 VDD.t1692 129.631
R1547 VDD.t1692 VDD.t201 129.631
R1548 VDD.t201 VDD.t1698 129.631
R1549 VDD.t1698 VDD.t189 129.631
R1550 VDD.t189 VDD.t1688 129.631
R1551 VDD.t1688 VDD.t4189 129.631
R1552 VDD.t4189 VDD.t2601 129.631
R1553 VDD.t2601 VDD.t4187 129.631
R1554 VDD.t4187 VDD.t1696 129.631
R1555 VDD.t1696 VDD.t4191 129.631
R1556 VDD.t4191 VDD.t1690 129.631
R1557 VDD.t1690 VDD.t4185 129.631
R1558 VDD.t4185 VDD.t1694 129.631
R1559 VDD.t3694 VDD.t1468 129.631
R1560 VDD.t2663 VDD.t2956 129.631
R1561 VDD.t3770 VDD.t3544 129.631
R1562 VDD.t1928 VDD.t3507 129.631
R1563 VDD.t3509 VDD.t1928 129.631
R1564 VDD.t1804 VDD.n1340 129.631
R1565 VDD.t3590 VDD.t856 129.631
R1566 VDD.t854 VDD.t3590 129.631
R1567 VDD.t394 VDD.t3776 129.631
R1568 VDD.t2759 VDD.t4294 129.631
R1569 VDD.t3578 VDD.t3206 129.631
R1570 VDD.t2780 VDD.t3045 129.631
R1571 VDD.t982 VDD.t3836 129.631
R1572 VDD.t1214 VDD.t3464 129.631
R1573 VDD.t2025 VDD.t1580 129.631
R1574 VDD.t4288 VDD.t2681 129.631
R1575 VDD.t2817 VDD.t3320 129.631
R1576 VDD.t2569 VDD.t3333 129.631
R1577 VDD.t2782 VDD.t2149 129.631
R1578 VDD.t2481 VDD.t1887 129.631
R1579 VDD.t2679 VDD.t3513 129.631
R1580 VDD.t1435 VDD.t2890 129.631
R1581 VDD.t3303 VDD.t3085 129.631
R1582 VDD.t1020 VDD.t941 129.631
R1583 VDD.t2151 VDD.t2249 129.631
R1584 VDD.t3747 VDD.t2182 129.631
R1585 VDD.t2129 VDD.t2391 129.631
R1586 VDD.t2363 VDD.t2134 129.631
R1587 VDD.t3821 VDD.t2888 129.631
R1588 VDD.t3915 VDD.t1986 129.631
R1589 VDD.t3846 VDD.t3202 129.631
R1590 VDD.t1500 VDD.t3531 129.631
R1591 VDD.t957 VDD.t3417 129.631
R1592 VDD.t2709 VDD.t3873 129.631
R1593 VDD.t3793 VDD.t3913 129.631
R1594 VDD.t2539 VDD.t2673 129.631
R1595 VDD.t1431 VDD.t2071 129.631
R1596 VDD.t2934 VDD.t1537 129.631
R1597 VDD.t2558 VDD.t1116 129.631
R1598 VDD.t701 VDD.t3390 129.631
R1599 VDD.t2999 VDD.t4022 129.631
R1600 VDD.t125 VDD.t43 129.631
R1601 VDD.t119 VDD.t117 129.631
R1602 VDD.t621 VDD.t41 129.631
R1603 VDD.t123 VDD.t121 129.631
R1604 VDD.t2608 VDD.t352 129.631
R1605 VDD.t2610 VDD.t319 129.631
R1606 VDD.t2634 VDD.t388 129.631
R1607 VDD.t2606 VDD.t354 129.631
R1608 VDD.t2614 VDD.t386 129.631
R1609 VDD.t2638 VDD.t347 129.631
R1610 VDD.t2612 VDD.t321 129.631
R1611 VDD.t2636 VDD.t390 129.631
R1612 VDD.t3789 VDD.t4290 129.631
R1613 VDD.t4211 VDD.t3173 129.631
R1614 VDD.t1473 VDD.t3246 129.631
R1615 VDD.t4266 VDD.t1354 129.631
R1616 VDD.t1207 VDD.t2013 129.631
R1617 VDD.t3250 VDD.t2483 129.631
R1618 VDD.t3132 VDD.t2395 129.631
R1619 VDD.n1175 VDD.t3764 129.631
R1620 VDD.t139 VDD.t1966 129.631
R1621 VDD.n1097 VDD.t4260 129.631
R1622 VDD.t1626 VDD.t2522 129.631
R1623 VDD.t2912 VDD.t2291 129.631
R1624 VDD.t2031 VDD.t2380 129.631
R1625 VDD.t1912 VDD.t3341 129.631
R1626 VDD.t1922 VDD.t3117 129.631
R1627 VDD.t3939 VDD.t3453 129.631
R1628 VDD.t1722 VDD.t1411 129.631
R1629 VDD.t1443 VDD.t2898 129.631
R1630 VDD.t1857 VDD.t4020 129.631
R1631 VDD.t2036 VDD.t1992 129.631
R1632 VDD.t4183 VDD.t1339 129.631
R1633 VDD.t4105 VDD.t2321 129.631
R1634 VDD.t4053 VDD.t2942 129.631
R1635 VDD.t1840 VDD.t3398 129.631
R1636 VDD.t3811 VDD.t3070 129.631
R1637 VDD.t2665 VDD.t2677 129.631
R1638 VDD.t2790 VDD.t3524 129.631
R1639 VDD.t2874 VDD.t3967 129.631
R1640 VDD.t4072 VDD.t3129 129.631
R1641 VDD.t1358 VDD.t2444 129.631
R1642 VDD.t2269 VDD.t1523 129.631
R1643 VDD.t1235 VDD.t3406 129.631
R1644 VDD.t4066 VDD.t2112 129.631
R1645 VDD.t3803 VDD.t4282 129.631
R1646 VDD.t2119 VDD.t3799 129.631
R1647 VDD.t2027 VDD.t1914 129.631
R1648 VDD.t3248 VDD.t4276 129.631
R1649 VDD.t2868 VDD.t998 129.631
R1650 VDD.t1291 VDD.t3567 129.631
R1651 VDD.t3576 VDD.t4040 129.631
R1652 VDD.t1865 VDD.t2330 129.631
R1653 VDD.t2675 VDD.t3007 129.631
R1654 VDD.t3154 VDD.t3682 129.631
R1655 VDD.t3515 VDD.t3108 129.631
R1656 VDD.t3353 VDD.t975 129.631
R1657 VDD.t1409 VDD.t2359 129.631
R1658 VDD.t2659 VDD.t3142 129.631
R1659 VDD.t3751 VDD.t4068 129.631
R1660 VDD.t2127 VDD.t3522 129.631
R1661 VDD.t2546 VDD.t2299 129.631
R1662 VDD.t3634 VDD.t3853 129.631
R1663 VDD.t3262 VDD.t1415 129.631
R1664 VDD.t3885 VDD.t1910 129.631
R1665 VDD.t4197 VDD.t1233 129.631
R1666 VDD.t3384 VDD.t2590 129.631
R1667 VDD.t2809 VDD.t3311 129.631
R1668 VDD.t2618 VDD.t3983 129.631
R1669 VDD.t3745 VDD.t2798 129.631
R1670 VDD.t2962 VDD.t1789 129.631
R1671 VDD.t2870 VDD.t2729 129.631
R1672 VDD.t1510 VDD.t2896 129.631
R1673 VDD.t2038 VDD.t2214 129.631
R1674 VDD.t3893 VDD.t2667 129.631
R1675 VDD.t1628 VDD.t977 129.631
R1676 VDD.t3198 VDD.t4038 129.631
R1677 VDD.t2361 VDD.t2368 129.631
R1678 VDD.t2669 VDD.t2251 129.631
R1679 VDD.t3949 VDD.t2253 129.631
R1680 VDD.t4042 VDD.t1682 129.631
R1681 VDD.t4096 VDD.t2860 129.631
R1682 VDD.t2489 VDD.t1231 129.631
R1683 VDD.t3686 VDD.t3279 129.631
R1684 VDD.t2493 VDD.t1800 129.631
R1685 VDD.t2757 VDD.t3574 129.631
R1686 VDD.t3572 VDD.t1812 129.631
R1687 VDD.t4199 VDD.t2101 129.631
R1688 VDD.t2277 VDD.t3087 129.631
R1689 VDD.t2450 VDD.t3986 129.631
R1690 VDD.t1718 VDD.t2807 129.631
R1691 VDD.t3586 VDD.t1810 129.631
R1692 VDD.t3591 VDD.t3419 129.631
R1693 VDD.t1134 VDD.t4207 129.631
R1694 VDD.t3074 VDD.t1481 129.631
R1695 VDD.t1582 VDD.t2800 129.631
R1696 VDD.t1138 VDD.t4201 129.631
R1697 VDD.t2725 VDD.t898 129.631
R1698 VDD.t3081 VDD.t4213 129.631
R1699 VDD.t1620 VDD.t3941 129.631
R1700 VDD.t3947 VDD.t3318 129.631
R1701 VDD.t2420 VDD.t2843 129.631
R1702 VDD.t1423 VDD.t1212 129.631
R1703 VDD.t1535 VDD.t3988 129.631
R1704 VDD.t1937 VDD.t1707 129.631
R1705 VDD.t3162 VDD.t3838 129.631
R1706 VDD.t2092 VDD.t3238 129.631
R1707 VDD.t2201 VDD.t2707 129.631
R1708 VDD.t3832 VDD.t4238 129.631
R1709 VDD.t1889 VDD.t2823 129.631
R1710 VDD.t3421 VDD.t2301 129.631
R1711 VDD.t2084 VDD.t3187 129.631
R1712 VDD.t4232 VDD.t3290 129.631
R1713 VDD.t984 VDD.t1730 129.631
R1714 VDD.t3684 VDD.t2835 129.631
R1715 VDD.t2029 VDD.t3457 129.631
R1716 VDD.t3369 VDD.t2061 129.631
R1717 VDD.t1984 VDD.t1777 129.631
R1718 VDD.t2554 VDD.t1479 129.631
R1719 VDD.t1739 VDD.t3049 129.631
R1720 VDD.t3640 VDD.t3469 129.631
R1721 VDD.t3923 VDD.t2157 129.631
R1722 VDD.t1259 VDD.t4177 129.631
R1723 VDD.t2560 VDD.t4171 129.631
R1724 VDD.t3665 VDD.t1226 129.631
R1725 VDD.t4227 VDD.t3112 129.631
R1726 VDD.t4167 VDD.t2125 129.631
R1727 VDD.t1245 VDD.t3381 129.631
R1728 VDD.t1228 VDD.t3688 129.631
R1729 VDD.t4011 VDD.t3536 129.631
R1730 VDD.t2642 VDD.t2721 129.631
R1731 VDD.t1297 VDD.t3451 129.631
R1732 VDD.t1251 VDD.t3345 129.631
R1733 VDD.t2172 VDD.t3091 129.631
R1734 VDD.t1370 VDD.t1679 129.631
R1735 VDD.t1195 VDD.t3976 129.631
R1736 VDD.t939 VDD.t965 129.631
R1737 VDD.t3528 VDD.t3929 129.631
R1738 VDD.t3377 VDD.t3999 129.631
R1739 VDD.t3252 VDD.t1732 129.631
R1740 VDD.t2640 VDD.t1737 129.631
R1741 VDD.t2520 VDD.t3136 129.631
R1742 VDD.t3714 VDD.t2434 129.631
R1743 VDD.t2829 VDD.t2007 129.631
R1744 VDD.t2661 VDD.t2209 129.631
R1745 VDD.t4286 VDD.t2159 129.631
R1746 VDD.t2902 VDD.t4280 129.631
R1747 VDD.t3102 VDD.t1099 129.631
R1748 VDD.t2398 VDD.t4076 129.631
R1749 VDD.t2303 VDD.t2448 129.631
R1750 VDD.t3881 VDD.t3236 129.631
R1751 VDD.t2839 VDD.t1632 129.631
R1752 VDD.t4101 VDD.t1684 129.631
R1753 VDD.t1982 VDD.t3842 129.631
R1754 VDD.t2954 VDD.t3003 129.631
R1755 VDD.t1350 VDD.t3277 129.631
R1756 VDD.t3005 VDD.t1802 129.631
R1757 VDD.t3425 VDD.t2900 129.631
R1758 VDD.t3152 VDD.t2476 129.631
R1759 VDD.t1990 VDD.t4218 129.631
R1760 VDD.t2042 VDD.t3654 129.631
R1761 VDD.t4169 VDD.t3718 129.631
R1762 VDD.t971 VDD.t2402 129.631
R1763 VDD.t3477 VDD.t2462 129.631
R1764 VDD.t4292 VDD.t3013 129.631
R1765 VDD.t4158 VDD.t1190 129.631
R1766 VDD.t2719 VDD.n2103 129.631
R1767 VDD.n2114 VDD.t1454 129.631
R1768 VDD.t3423 VDD.t3449 129.631
R1769 VDD.t1332 VDD.t3805 129.631
R1770 VDD.t3963 VDD.t3642 129.631
R1771 VDD.t1616 VDD.t4163 129.631
R1772 VDD.t3995 VDD.t4156 129.631
R1773 VDD.t3041 VDD.t1224 129.631
R1774 VDD.t4225 VDD.t3110 129.631
R1775 VDD.t4150 VDD.t2275 129.631
R1776 VDD.t1097 VDD.t1761 129.631
R1777 VDD.t1417 VDD.t1289 129.631
R1778 VDD.t1832 VDD.t2944 129.631
R1779 VDD.t2372 VDD.t2297 129.631
R1780 VDD.t933 VDD.t3178 129.631
R1781 VDD.t1247 VDD.t3636 129.631
R1782 VDD.t2063 VDD.t1179 129.631
R1783 VDD.t2652 VDD.t1249 129.631
R1784 VDD.t1421 VDD.t2207 129.631
R1785 VDD.t2485 VDD.t1388 129.631
R1786 VDD.t2991 VDD.t1674 129.631
R1787 VDD.t3971 VDD.t3373 129.631
R1788 VDD.t1724 VDD.t2703 129.631
R1789 VDD.t3427 VDD.t2603 129.631
R1790 VDD.t2872 VDD.t2422 129.631
R1791 VDD.t2533 VDD.t4103 129.631
R1792 VDD.t1975 VDD.t3158 129.631
R1793 VDD.t3455 VDD.t3671 129.631
R1794 VDD.t1433 VDD.t2575 129.631
R1795 VDD.t3404 VDD.t3435 129.631
R1796 VDD.t2537 VDD.t3266 129.631
R1797 VDD.t3484 VDD.t3584 129.631
R1798 VDD.t3787 VDD.t3034 129.631
R1799 VDD.t914 VDD.t1241 129.631
R1800 VDD.t3240 VDD.t3809 129.631
R1801 VDD.t2815 VDD.t923 129.631
R1802 VDD.t3100 VDD.t3937 129.631
R1803 VDD.t4203 VDD.t3379 129.631
R1804 VDD.t959 VDD.t3679 129.631
R1805 VDD.t1769 VDD.t3269 129.631
R1806 VDD.t1471 VDD.t2864 129.631
R1807 VDD.t4270 VDD.t1345 129.631
R1808 VDD.t2831 VDD.t1900 129.631
R1809 VDD.t1557 VDD.t4005 129.631
R1810 VDD.t3119 VDD.t3673 129.631
R1811 VDD.t3371 VDD.t2821 129.631
R1812 VDD.t1186 VDD.t1321 129.631
R1813 VDD.t2849 VDD.t3867 129.631
R1814 VDD.t2414 VDD.t2958 129.631
R1815 VDD.t3712 VDD.t918 129.631
R1816 VDD.t935 VDD.t927 129.631
R1817 VDD.t1498 VDD.t2979 129.631
R1818 VDD.t3441 VDD.t1343 129.631
R1819 VDD.t3593 VDD.t2579 129.631
R1820 VDD.t1136 VDD.t3917 129.631
R1821 VDD.t1979 VDD.t2404 129.631
R1822 VDD.t1539 VDD.t2833 129.631
R1823 VDD.t2216 VDD.t2966 129.631
R1824 VDD.t3160 VDD.t4143 129.631
R1825 VDD.t2845 VDD.t1149 129.631
R1826 VDD.t3164 VDD.t3367 129.631
R1827 VDD.t1437 VDD.t2491 129.631
R1828 VDD.t1793 VDD.t3935 129.631
R1829 VDD.t3830 VDD.t2894 129.631
R1830 VDD.t3305 VDD.t3827 129.631
R1831 VDD.t904 VDD.t1945 129.631
R1832 VDD.t3778 VDD.t1634 129.631
R1833 VDD.t3877 VDD.t3166 129.631
R1834 VDD.t874 VDD.t1898 129.631
R1835 VDD.t3171 VDD.t1280 129.631
R1836 VDD.t2516 VDD.t1103 129.631
R1837 VDD.t2271 VDD.t2468 129.631
R1838 VDD.t2203 VDD.t1105 129.631
R1839 VDD.t2153 VDD.t3314 129.631
R1840 VDD.t2090 VDD.t3180 129.631
R1841 VDD.t2220 VDD.t1575 129.631
R1842 VDD.t2273 VDD.t2472 129.631
R1843 VDD.t2264 VDD.t3169 129.631
R1844 VDD.t2571 VDD.t3146 129.631
R1845 VDD.t1988 VDD.t1142 129.631
R1846 VDD.t1969 VDD.t2174 129.631
R1847 VDD.n651 VDD.t4048 129.631
R1848 VDD.t900 VDD.n652 129.631
R1849 VDD.n653 VDD.t4015 129.631
R1850 VDD.n219 VDD.t2046 129.631
R1851 VDD.t2236 VDD.n218 129.631
R1852 VDD.t1401 VDD.n2277 129.631
R1853 VDD.n2278 VDD.t4003 129.631
R1854 VDD.t4055 VDD.n2279 129.631
R1855 VDD.t4001 VDD.t3351 129.631
R1856 VDD.n2281 VDD.t2196 129.631
R1857 VDD.t2074 VDD.t2505 128.472
R1858 VDD.t1427 VDD.t726 128.472
R1859 VDD.t1396 VDD.t3121 128.472
R1860 VDD.t3675 VDD.t2212 128.472
R1861 VDD.t461 VDD.t3232 128.472
R1862 VDD.t637 VDD.t3580 127.316
R1863 VDD.t1548 VDD.t4063 127.316
R1864 VDD.t3309 VDD.t471 127.316
R1865 VDD.t479 VDD.t3479 126.157
R1866 VDD.t706 VDD.t2723 126.157
R1867 VDD.t466 VDD.t511 126.157
R1868 VDD.t1906 VDD.t860 125.15
R1869 VDD.t756 VDD.t17 125.001
R1870 VDD.t571 VDD.t1109 125.001
R1871 VDD.t3196 VDD.t1270 123.844
R1872 VDD.t3616 VDD.t2535 123.844
R1873 VDD.t3389 VDD.t3337 123.844
R1874 VDD.t1336 VDD.t3760 123.844
R1875 VDD.t1334 VDD.t3761 123.844
R1876 VDD.t2246 VDD.t3758 123.844
R1877 VDD.t787 VDD.t351 123.844
R1878 VDD.t4092 VDD.n409 122.686
R1879 VDD.t1428 VDD.t892 121.528
R1880 VDD.t3031 VDD.t3054 121.528
R1881 VDD.t1485 VDD.t2743 121.528
R1882 VDD.t3598 VDD.t719 121.528
R1883 VDD.t2746 VDD.t3061 120.371
R1884 VDD.t1347 VDD.t3444 120.371
R1885 VDD.t1463 VDD.t1203 120.371
R1886 VDD.t1382 VDD.t1784 119.475
R1887 VDD.t527 VDD.t1266 119.213
R1888 VDD.t1025 VDD.t1830 118.281
R1889 VDD.t3669 VDD.t4070 118.281
R1890 VDD.t3696 VDD.t362 118.056
R1891 VDD.t1468 VDD.t3696 118.056
R1892 VDD.t4014 VDD.t3051 118.056
R1893 VDD.t1157 VDD.t3244 118.056
R1894 VDD.t2145 VDD.t2655 118.056
R1895 VDD.t4244 VDD.t1265 118.056
R1896 VDD.t1603 VDD.t929 116.898
R1897 VDD.t1670 VDD.t1880 116.898
R1898 VDD.t3743 VDD.t3849 116.898
R1899 VDD.t534 VDD.t1578 116.898
R1900 VDD.t3490 VDD.t3503 116.898
R1901 VDD.t3061 VDD.t3879 115.742
R1902 VDD.t862 VDD.t1599 115.742
R1903 VDD.t1490 VDD.t71 115.742
R1904 VDD.t4274 VDD.t63 115.742
R1905 VDD.t751 VDD.t287 115.742
R1906 VDD.t3952 VDD.t3489 115.742
R1907 VDD.t413 VDD.t649 115.742
R1908 VDD.t3364 VDD.t311 115.742
R1909 VDD.t2138 VDD.t1873 115.742
R1910 VDD.t892 VDD.t3965 114.584
R1911 VDD.t3054 VDD.t3801 114.584
R1912 VDD.t360 VDD.t1485 114.584
R1913 VDD.t3517 VDD.n325 114.584
R1914 VDD.t719 VDD.t15 114.584
R1915 VDD.t1164 VDD.t2355 114.422
R1916 VDD.n494 VDD.t2803 113.427
R1917 VDD.t4082 VDD.n409 113.427
R1918 VDD.t4173 VDD.t1554 113.427
R1919 VDD.t3329 VDD.t2859 113.427
R1920 VDD.t1676 VDD.t1323 113.209
R1921 VDD.t1122 VDD.t3648 112.269
R1922 VDD.t3337 VDD.t3616 112.269
R1923 VDD.t2706 VDD.t3389 112.269
R1924 VDD.t351 VDD.t2562 112.269
R1925 VDD.t2142 VDD.t1836 112.269
R1926 VDD.t646 VDD.t2595 111.112
R1927 VDD.t2241 VDD.t1193 111.112
R1928 VDD.t1272 VDD.t1954 109.954
R1929 VDD.t1274 VDD.t605 109.954
R1930 VDD.t2503 VDD.t466 109.954
R1931 VDD.t440 VDD.t637 108.796
R1932 VDD.t4063 VDD.t0 108.796
R1933 VDD.t471 VDD.t1453 108.796
R1934 VDD.t1392 VDD.t1767 107.639
R1935 VDD.t2713 VDD.t356 106.481
R1936 VDD.t191 VDD.t1943 106.481
R1937 VDD.t1656 VDD.t2974 106.481
R1938 VDD.t2742 VDD.t3509 106.481
R1939 VDD.t3866 VDD.t854 106.481
R1940 VDD.t3776 VDD.t2356 106.481
R1941 VDD.t1614 VDD.t3632 106.481
R1942 VDD.t3394 VDD.t701 106.481
R1943 VDD.t41 VDD.t119 106.481
R1944 VDD.t388 VDD.t2610 106.481
R1945 VDD.t386 VDD.t2606 106.481
R1946 VDD.t321 VDD.t2638 106.481
R1947 VDD.t790 VDD.t1774 106.481
R1948 VDD.t3983 VDD.t3475 106.481
R1949 VDD.t2035 VDD.t3714 106.481
R1950 VDD.t3446 VDD.t1853 105.325
R1951 VDD.t3429 VDD.t1927 105.325
R1952 VDD.t3871 VDD.t2438 105.325
R1953 VDD.t3499 VDD.t1517 105.325
R1954 VDD.t1568 VDD.t434 105.138
R1955 VDD.t906 VDD.t2225 105.138
R1956 VDD.t4175 VDD.t3973 104.168
R1957 VDD.t758 VDD.t443 104.168
R1958 VDD.t3150 VDD.t2685 104.168
R1959 VDD.t1111 VDD.t3907 103.01
R1960 VDD.t2382 VDD.n1857 103.01
R1961 VDD.t1276 VDD.t3582 103.01
R1962 VDD.t3957 VDD.t1601 101.853
R1963 VDD.t3834 VDD.t3710 101.853
R1964 VDD.t2358 VDD.t1614 101.853
R1965 VDD.t773 VDD.t279 101.853
R1966 VDD.t2474 VDD.t1465 101.853
R1967 VDD.t3690 VDD.t2588 101.853
R1968 VDD.t2593 VDD.t1885 100.695
R1969 VDD.t2592 VDD.t1884 100.695
R1970 VDD.t636 VDD.t1512 100.695
R1971 VDD.t4035 VDD.t467 99.5375
R1972 VDD.t979 VDD.t2454 99.5375
R1973 VDD.t323 VDD.t3772 99.5375
R1974 VDD.t537 VDD.n1669 98.9278
R1975 VDD.t3720 VDD.t1230 98.3801
R1976 VDD.t3823 VDD.t1870 98.3801
R1977 VDD.t3731 VDD.t3757 98.3801
R1978 VDD.t2076 VDD.t3106 98.3801
R1979 VDD.t1783 VDD.t1384 97.2227
R1980 VDD.t689 VDD.t2121 97.2227
R1981 VDD.t648 VDD.t4195 97.2227
R1982 VDD.t3079 VDD.t1950 96.0653
R1983 VDD.t185 VDD.t3094 96.0653
R1984 VDD.t1077 VDD.t800 95.3521
R1985 VDD.t2452 VDD.t979 94.9079
R1986 VDD.t2454 VDD.t980 94.9079
R1987 VDD.t3534 VDD.t2295 94.9079
R1988 VDD.t3386 VDD.t3701 94.9079
R1989 VDD.t1884 VDD.t2593 93.7505
R1990 VDD.t1664 VDD.t994 93.7505
R1991 VDD.t3741 VDD.t1569 93.7505
R1992 VDD.t3768 VDD.t449 92.5931
R1993 VDD.t392 VDD.t1586 92.5931
R1994 VDD.t613 VDD.t4133 92.5931
R1995 VDD.t26 VDD.t807 92.5931
R1996 VDD.t1086 VDD.t813 92.5931
R1997 VDD.t1060 VDD.t597 92.5931
R1998 VDD.t1058 VDD.t1088 92.5931
R1999 VDD.t1090 VDD.t2050 92.5931
R2000 VDD.t825 VDD.t4127 92.5931
R2001 VDD.t3299 VDD.t4118 92.5931
R2002 VDD.t2626 VDD.t416 92.5931
R2003 VDD.t2630 VDD.t305 92.5931
R2004 VDD.t2587 VDD.t3690 92.5931
R2005 VDD.t2628 VDD.t2005 92.5931
R2006 VDD.t3612 VDD.t3990 92.5931
R2007 VDD.t3652 VDD.t1513 90.801
R2008 VDD.t3089 VDD.t4179 90.801
R2009 VDD.t747 VDD.t732 90.2783
R2010 VDD.n1272 VDD.t3023 90.2783
R2011 VDD.t3388 VDD.t1044 90.2783
R2012 VDD.t4260 VDD.t2528 90.2783
R2013 VDD.t3975 VDD.t4175 90.2783
R2014 VDD.t1715 VDD.t925 89.6062
R2015 VDD.t1925 VDD.t3429 89.1209
R2016 VDD.t633 VDD.t1326 89.1209
R2017 VDD.t203 VDD.t1486 87.9635
R2018 VDD.t1686 VDD.t2768 87.9635
R2019 VDD.t3632 VDD.t1613 87.9635
R2020 VDD.t2244 VDD.t2238 87.9635
R2021 VDD.t1676 VDD.n2109 87.1921
R2022 VDD.t4216 VDD.t3980 86.8061
R2023 VDD.t2936 VDD.t741 85.6486
R2024 VDD.t4258 VDD.t1960 85.6486
R2025 VDD.t1413 VDD.t2727 85.6486
R2026 VDD.t3375 VDD.t1700 84.4912
R2027 VDD.t767 VDD.t4024 84.4912
R2028 VDD.t3659 VDD.t861 84.4912
R2029 VDD.t1953 VDD.t1272 84.4912
R2030 VDD.t3498 VDD.t463 84.4912
R2031 VDD.t3755 VDD.t445 84.4912
R2032 VDD.t324 VDD.t3610 83.3338
R2033 VDD.t703 VDD.t4033 83.3338
R2034 VDD.t1222 VDD.t638 83.3338
R2035 VDD.t2753 VDD.t4117 83.3338
R2036 VDD.t3 VDD.t1132 83.3338
R2037 VDD.t2057 VDD.t4240 83.3338
R2038 VDD.t4139 VDD.t496 83.3338
R2039 VDD.t4062 VDD.t1441 83.3338
R2040 VDD.t3546 VDD.t2226 82.1764
R2041 VDD.t426 VDD.t3921 81.243
R2042 VDD.t2857 VDD.t3329 81.019
R2043 VDD.t3965 VDD.t890 79.8616
R2044 VDD.n610 VDD.t736 79.8616
R2045 VDD.t4250 VDD.n510 79.8616
R2046 VDD.t1605 VDD.t3322 79.8616
R2047 VDD.t792 VDD.t2117 79.8616
R2048 VDD.t3749 VDD.t2847 79.8616
R2049 VDD.t1380 VDD.t763 78.7042
R2050 VDD.t1255 VDD.t293 78.7042
R2051 VDD.t4261 VDD.t285 78.7042
R2052 VDD.t418 VDD.t3307 77.5468
R2053 VDD.t4120 VDD.t4046 77.5468
R2054 VDD.t1577 VDD.t534 77.5468
R2055 VDD.t3244 VDD.t1155 76.3894
R2056 VDD.t2655 VDD.t2144 76.3894
R2057 VDD.t2654 VDD.t2145 76.3894
R2058 VDD.t2524 VDD.t1168 75.232
R2059 VDD.t1531 VDD.t24 75.232
R2060 VDD.t2293 VDD.t447 74.0746
R2061 VDD.t4018 VDD.t1378 74.0746
R2062 VDD.t1592 VDD.t1563 74.0746
R2063 VDD.t615 VDD.t1446 74.0746
R2064 VDD.t4147 VDD.t2168 74.0746
R2065 VDD.t2788 VDD.t3360 74.0746
R2066 VDD.t155 VDD.t2507 74.0746
R2067 VDD.t3840 VDD.t28 74.0746
R2068 VDD.t817 VDD.t2882 74.0746
R2069 VDD.t177 VDD.t153 74.0746
R2070 VDD.t171 VDD.t149 74.0746
R2071 VDD.t3064 VDD.t3630 74.0746
R2072 VDD.t486 VDD.t1867 74.0746
R2073 VDD.n601 VDD.t13 72.9172
R2074 VDD.t3053 VDD.t3031 72.9172
R2075 VDD.t2743 VDD.t1483 72.9172
R2076 VDD.t3230 VDD.t3316 72.9172
R2077 VDD.t181 VDD.t1036 72.9172
R2078 VDD.t1072 VDD.t1470 72.8798
R2079 VDD.t53 VDD.t1824 71.7598
R2080 VDD.t2495 VDD.t2581 71.7598
R2081 VDD.t2892 VDD.t4036 71.7598
R2082 VDD.t1451 VDD.t1996 71.7598
R2083 VDD.t2573 VDD.t1814 71.7598
R2084 VDD.t1269 VDD.t3196 70.6024
R2085 VDD.t3729 VDD.t3862 70.6024
R2086 VDD.t601 VDD.t1068 70.6024
R2087 VDD.t3761 VDD.t1336 70.6024
R2088 VDD.t3622 VDD.t3338 70.4903
R2089 VDD.t1776 VDD.t1430 69.4449
R2090 VDD.t318 VDD.t1467 69.4449
R2091 VDD.t603 VDD.t2904 69.4449
R2092 VDD.t821 VDD.t1166 69.4449
R2093 VDD.t1295 VDD.t916 69.4449
R2094 VDD.t2632 VDD.t2740 69.4449
R2095 VDD.t3825 VDD.t4284 69.4449
R2096 VDD.t2082 VDD.t2854 69.4449
R2097 VDD.t3123 VDD.t4193 69.4449
R2098 VDD.t1977 VDD.t631 68.1009
R2099 VDD.t809 VDD.t780 67.7513
R2100 VDD.t3281 VDD.t1826 67.1301
R2101 VDD.t3283 VDD.t1828 67.1301
R2102 VDD.t2319 VDD.t1349 67.1301
R2103 VDD.t2083 VDD.n303 67.1301
R2104 VDD.t1962 VDD.t2461 67.1301
R2105 VDD.n255 VDD.t3991 67.1301
R2106 VDD.t3905 VDD.t3560 66.9061
R2107 VDD.t1720 VDD.t1386 66.9061
R2108 VDD.t2671 VDD.t945 66.9061
R2109 VDD.t3339 VDD.t1971 66.9061
R2110 VDD.t2505 VDD.t2073 65.9727
R2111 VDD.t2408 VDD.t1074 65.9727
R2112 VDD.t3121 VDD.t1395 65.9727
R2113 VDD.t1822 VDD.t1199 65.9727
R2114 VDD.t3505 VDD.t798 65.7114
R2115 VDD.t2332 VDD.t3628 64.8153
R2116 VDD.t754 VDD.t420 64.8153
R2117 VDD.t531 VDD.t1495 64.8153
R2118 VDD.t1171 VDD.t477 64.8153
R2119 VDD.t309 VDD.t517 64.8153
R2120 VDD.t1920 VDD.t497 64.8153
R2121 VDD.t1705 VDD.t1366 63.6579
R2122 VDD.t4007 VDD.t2866 63.6579
R2123 VDD.t2805 VDD.t519 62.5005
R2124 VDD.t1267 VDD.t3182 62.5005
R2125 VDD.t644 VDD.t2556 62.5005
R2126 VDD.t2564 VDD.t3597 62.5005
R2127 VDD.t525 VDD.t1837 62.5005
R2128 VDD.n621 VDD.t57 62.1822
R2129 VDD.t2964 VDD.t30 62.1271
R2130 VDD.t1931 VDD.n350 62.1271
R2131 VDD.t4026 VDD.t1040 61.979
R2132 VDD.t1325 VDD.t2015 61.3431
R2133 VDD.t2827 VDD.t536 61.3431
R2134 VDD.t2478 VDD.t1728 60.9324
R2135 VDD.t2430 VDD.t3437 60.1857
R2136 VDD.t743 VDD.t1390 60.1857
R2137 VDD.t3753 VDD.t1672 60.1857
R2138 VDD.t2442 VDD.t2649 59.0283
R2139 VDD.t3782 VDD.n1598 59.0283
R2140 VDD.t878 VDD.t3705 59.0283
R2141 VDD.t877 VDD.t3703 59.0283
R2142 VDD.n577 VDD.t1124 57.8709
R2143 VDD.n600 VDD.t199 57.8709
R2144 VDD.t1566 VDD.n586 57.8709
R2145 VDD.t1816 VDD.n401 57.8709
R2146 VDD.n1775 VDD.t611 57.8709
R2147 VDD.t3487 VDD.t1184 57.8709
R2148 VDD.t2997 VDD.t2416 57.8709
R2149 VDD.t4107 VDD.t1881 57.8709
R2150 VDD.t3558 VDD.t2233 57.8709
R2151 VDD.t2400 VDD.t4242 57.8709
R2152 VDD.t4268 VDD.t4246 57.8709
R2153 VDD.t1933 VDD.t1012 57.8709
R2154 VDD.t2884 VDD.t1004 57.8709
R2155 VDD.t4051 VDD.t1018 57.8709
R2156 VDD.t1662 VDD.t1008 57.8709
R2157 VDD.t1205 VDD.t888 57.8709
R2158 VDD.t3226 VDD.t884 57.8709
R2159 VDD.t2938 VDD.t655 57.8709
R2160 VDD.t1851 VDD.t623 57.8709
R2161 VDD.t4099 VDD.t665 57.8709
R2162 VDD.t3774 VDD.t627 57.8709
R2163 VDD.t2104 VDD.t2984 56.7135
R2164 VDD.t1064 VDD.t1861 56.7135
R2165 VDD.t2163 VDD.t1999 56.7135
R2166 VDD.t3600 VDD.t2543 56.7135
R2167 VDD.t1908 VDD.t503 56.7135
R2168 VDD.t3903 VDD.t902 55.5561
R2169 VDD.t3218 VDD.t3287 55.5561
R2170 VDD.t2541 VDD.t3443 55.5561
R2171 VDD.t852 VDD.t3993 55.5561
R2172 VDD.t2705 VDD.t3624 55.5561
R2173 VDD.t143 VDD.t1968 55.5561
R2174 VDD.t3096 VDD.t1033 55.5561
R2175 VDD.t575 VDD.t1869 54.3986
R2176 VDD.t1712 VDD.t1181 53.2412
R2177 VDD.t1493 VDD.t1177 52.5692
R2178 VDD.t1093 VDD.t1666 52.5692
R2179 VDD.t3791 VDD.t3739 52.5692
R2180 VDD.t3447 VDD.t1855 52.0838
R2181 VDD.t4028 VDD.t2328 52.0838
R2182 VDD.t783 VDD.t3780 52.0838
R2183 VDD.t708 VDD.t3897 50.9264
R2184 VDD.t3663 VDD.t1895 50.9264
R2185 VDD.t3220 VDD.t3260 50.9264
R2186 VDD.t2993 VDD.t4084 50.9264
R2187 VDD.t2326 VDD.t4080 50.9264
R2188 VDD.t4086 VDD.t335 50.9264
R2189 VDD.t187 VDD.t147 50.9264
R2190 VDD.t175 VDD.t145 50.9264
R2191 VDD.t2879 VDD.t2886 50.9264
R2192 VDD.t2928 VDD.t1113 50.9264
R2193 VDD.t1095 VDD.t2922 50.9264
R2194 VDD.t2170 VDD.t2733 49.769
R2195 VDD.t2240 VDD.t2970 48.985
R2196 VDD.t1894 VDD.n525 48.8682
R2197 VDD.t710 VDD.t1031 48.6116
R2198 VDD.t2851 VDD.t1399 47.4542
R2199 VDD.t1042 VDD.t617 46.9764
R2200 VDD.t3293 VDD.t3795 46.2968
R2201 VDD.t3727 VDD.t3224 46.2968
R2202 VDD.t609 VDD.t3393 46.2968
R2203 VDD.t480 VDD.t1243 46.2968
R2204 VDD.t4121 VDD.t2393 46.2968
R2205 VDD.t4064 VDD.t3015 46.2968
R2206 VDD.t1054 VDD.t642 46.2968
R2207 VDD.t469 VDD.t1261 45.1394
R2208 VDD.t2986 VDD.t717 43.982
R2209 VDD.t948 VDD.t3285 43.982
R2210 VDD.n334 VDD.t1916 43.982
R2211 VDD.t4257 VDD.t2624 43.982
R2212 VDD.t3234 VDD.n473 42.8246
R2213 VDD.t523 VDD.t663 42.8246
R2214 VDD.t802 VDD.t804 41.6672
R2215 VDD.t1716 VDD.t2065 41.6672
R2216 VDD.t475 VDD.t3242 41.6672
R2217 VDD.t2136 VDD.t83 41.6672
R2218 VDD.t297 VDD.t283 41.6672
R2219 VDD.t291 VDD.t1284 41.6672
R2220 VDD.t3860 VDD.t4209 41.6672
R2221 VDD.t1120 VDD.t303 41.6672
R2222 VDD.t2432 VDD.t3077 41.6672
R2223 VDD.t1506 VDD.t236 41.6672
R2224 VDD.t3850 VDD.t2003 41.6672
R2225 VDD.t490 VDD.t2231 41.6672
R2226 VDD.t2737 VDD.t1640 41.6672
R2227 VDD.t2734 VDD.t1644 41.6672
R2228 VDD.t3431 VDD.n566 40.5098
R2229 VDD.t3602 VDD.n576 40.5098
R2230 VDD.t2972 VDD.t2262 40.5098
R2231 VDD.n1265 VDD.t1151 40.5098
R2232 VDD.t3961 VDD.n1776 40.5098
R2233 VDD.t3030 VDD.t1711 38.1949
R2234 VDD.t1807 VDD.t695 38.1949
R2235 VDD.t3959 VDD.t659 38.1949
R2236 VDD.t2334 VDD.t2184 37.0375
R2237 VDD.t1652 VDD.t4123 37.0375
R2238 VDD.t858 VDD.t1263 37.0375
R2239 VDD.t4205 VDD.t2189 37.0375
R2240 VDD.t3486 VDD.t2616 37.0375
R2241 VDD.t1192 VDD.t2188 37.0375
R2242 VDD.t1504 VDD.t2550 37.0375
R2243 VDD.t775 VDD.t1959 37.0375
R2244 VDD.t3646 VDD.t432 35.8801
R2245 VDD.t3019 VDD.t2052 35.8801
R2246 VDD.t2466 VDD.t1211 34.7227
R2247 VDD.t2968 VDD.t1140 34.7227
R2248 VDD.t4078 VDD.t281 34.7227
R2249 VDD.t2622 VDD.t1791 34.7227
R2250 VDD.t1779 VDD.t3618 34.6481
R2251 VDD.t1253 VDD.t3402 33.5653
R2252 VDD.t3657 VDD.t2908 33.5653
R2253 VDD.t3362 VDD.t2198 33.5653
R2254 VDD.t749 VDD.t973 33.5653
R2255 VDD.t3895 VDD.t2512 32.4079
R2256 VDD.t2566 VDD.t3039 32.4079
R2257 VDD.t165 VDD.t829 32.4079
R2258 VDD.t163 VDD.t827 32.4079
R2259 VDD.t159 VDD.t837 32.4079
R2260 VDD.t161 VDD.t841 32.4079
R2261 VDD.t1286 VDD.t295 32.4079
R2262 VDD.t2751 VDD.t299 32.4079
R2263 VDD.t3474 VDD.t410 32.4079
R2264 VDD.t3583 VDD.t439 32.4079
R2265 VDD.t3887 VDD.t3177 32.4079
R2266 VDD.t1000 VDD.t1126 31.2505
R2267 VDD.t2499 VDD.t3415 31.2505
R2268 VDD.t3114 VDD.t1081 31.2505
R2269 VDD.t2914 VDD.t1702 31.2505
R2270 VDD.t3254 VDD.t4114 31.2505
R2271 VDD.t746 VDD.t2748 31.2505
R2272 VDD.t4154 VDD.t3466 31.2505
R2273 VDD.t3347 VDD.t3140 30.0931
R2274 VDD.t3026 VDD.t725 30.0931
R2275 VDD.t1183 VDD.t3275 30.0931
R2276 VDD.t1544 VDD.t2976 28.9357
R2277 VDD.t3588 VDD.t3501 28.9357
R2278 VDD.t2745 VDD.t1101 28.6743
R2279 VDD.t661 VDD.t1965 28.6743
R2280 VDD.t1175 VDD.t1489 28.6743
R2281 VDD.t1668 VDD.t3363 28.6743
R2282 VDD.t3737 VDD.t2140 28.6743
R2283 VDD.t1941 VDD.t713 27.7783
R2284 VDD.t2518 VDD.t3265 27.7783
R2285 VDD.t69 VDD.t910 27.7783
R2286 VDD.t315 VDD.t2176 27.7783
R2287 VDD.t2059 VDD.t2853 27.7783
R2288 VDD.t1877 VDD.t1533 27.7783
R2289 VDD.t1323 VDD.n2115 27.4448
R2290 VDD.t1376 VDD.t2747 26.6209
R2291 VDD.t2186 VDD.t3033 26.6209
R2292 VDD.t4222 VDD.t1973 26.6209
R2293 VDD.t4109 VDD.t4060 26.6209
R2294 VDD.t522 VDD.t9 26.6209
R2295 VDD.t2 VDD.t1362 25.4635
R2296 VDD.t1356 VDD.t2459 25.4635
R2297 VDD.t786 VDD.n348 25.0303
R2298 VDD.t4125 VDD.t3057 23.1486
R2299 VDD.t5 VDD.t1588 23.1486
R2300 VDD.t437 VDD.t1590 23.1486
R2301 VDD.t3358 VDD.t1107 23.1486
R2302 VDD.t1552 VDD.t805 23.1486
R2303 VDD.t759 VDD.t2819 23.1486
R2304 VDD.t645 VDD.t2620 23.1486
R2305 VDD.n262 VDD.t2683 21.9912
R2306 VDD.t727 VDD.t1556 20.8338
R2307 VDD.t1735 VDD.t3570 20.8338
R2308 VDD.t1734 VDD.t3569 20.8338
R2309 VDD.t1543 VDD.t1947 20.8338
R2310 VDD.t1541 VDD.t1948 20.8338
R2311 VDD.n348 VDD.t955 19.2958
R2312 VDD.n350 VDD.t996 18.8763
R2313 VDD.t3214 VDD.t4131 18.519
R2314 VDD.t3331 VDD.t4141 18.519
R2315 VDD.t1714 VDD.t3488 18.519
R2316 VDD.t1492 VDD.t67 18.519
R2317 VDD.n1098 VDD.n1097 18.519
R2318 VDD.t3366 VDD.t301 18.519
R2319 VDD.t2141 VDD.t2001 18.519
R2320 VDD.t2374 VDD.n342 16.7667
R2321 VDD.t1330 VDD.t3295 16.2042
R2322 VDD.t2103 VDD.t4129 15.0468
R2323 VDD.t515 VDD.t4224 15.0468
R2324 VDD.t442 VDD.t509 15.0468
R2325 VDD.t2406 VDD.t2916 15.0468
R2326 VDD.t844 VDD.t499 15.0468
R2327 VDD.t1257 VDD.t3194 15.0468
R2328 VDD.t2513 VDD.t3899 14.3374
R2329 VDD.t1278 VDD.t1497 14.3374
R2330 VDD.t504 VDD.t3481 14.3032
R2331 VDD.t1611 VDD.t2711 13.8894
R2332 VDD.t699 VDD.t481 13.8894
R2333 VDD.n919 VDD.t3184 13.8894
R2334 VDD.n1607 VDD.t1957 12.8338
R2335 VDD.n437 VDD.t1400 12.8338
R2336 VDD.n338 VDD.t3131 12.8338
R2337 VDD.n918 VDD.t2858 12.8338
R2338 VDD.n266 VDD.t1210 12.8338
R2339 VDD.t3958 VDD.t424 12.732
R2340 VDD.t3891 VDD.t4234 12.732
R2341 VDD.t3047 VDD.t1279 12.732
R2342 VDD.t539 VDD.t3750 12.732
R2343 VDD.n544 VDD.n527 11.8275
R2344 VDD.n1662 VDD.n467 11.8275
R2345 VDD.n564 VDD.t3668 11.8234
R2346 VDD.n1375 VDD.t2261 11.8234
R2347 VDD.n1390 VDD.t2162 11.8234
R2348 VDD.n504 VDD.t419 11.8234
R2349 VDD.n511 VDD.t1768 11.8234
R2350 VDD.n515 VDD.t3084 11.8234
R2351 VDD.n1389 VDD.t4221 11.8234
R2352 VDD.n1345 VDD.t2578 11.8234
R2353 VDD.n1351 VDD.t3872 11.8234
R2354 VDD.n492 VDD.t2863 11.8234
R2355 VDD.n1600 VDD.t2118 11.8234
R2356 VDD.n1609 VDD.t2789 11.8234
R2357 VDD.n1601 VDD.t2390 11.8234
R2358 VDD.n485 VDD.t2329 11.8234
R2359 VDD.n490 VDD.t2320 11.8234
R2360 VDD.n1264 VDD.t1450 11.8234
R2361 VDD.n468 VDD.t4235 11.8234
R2362 VDD.n438 VDD.t2852 11.8234
R2363 VDD.n435 VDD.t3845 11.8234
R2364 VDD.n1177 VDD.t1200 11.8234
R2365 VDD.n1791 VDD.t1831 11.8234
R2366 VDD.n371 VDD.t2887 11.8234
R2367 VDD.n370 VDD.t2929 11.8234
R2368 VDD.n377 VDD.t881 11.8234
R2369 VDD.n324 VDD.t1119 11.8234
R2370 VDD.n339 VDD.t1445 11.8234
R2371 VDD.n345 VDD.t4071 11.8234
R2372 VDD.n336 VDD.t2375 11.8234
R2373 VDD.n328 VDD.t3956 11.8234
R2374 VDD.n1954 VDD.t2437 11.8234
R2375 VDD.n1953 VDD.t3596 11.8234
R2376 VDD.n916 VDD.t3535 11.8234
R2377 VDD.n301 VDD.t2551 11.8234
R2378 VDD.n294 VDD.t3233 11.8234
R2379 VDD.n922 VDD.t3356 11.8234
R2380 VDD.n265 VDD.t2232 11.8234
R2381 VDD.n258 VDD.t3613 11.8234
R2382 VDD.n2107 VDD.t2245 11.8234
R2383 VDD.t3462 VDD.t753 11.5746
R2384 VDD.t1676 VDD.n2114 11.5746
R2385 VDD.t2464 VDD.t641 11.5746
R2386 VDD.t472 VDD.t349 11.5746
R2387 VDD.n1527 VDD.t734 11.0764
R2388 VDD.n1663 VDD.t505 11.0764
R2389 VDD.t1930 VDD.t786 10.6968
R2390 VDD.t3608 VDD.t778 10.4172
R2391 VDD.t2376 VDD.t1935 10.4172
R2392 VDD.t3526 VDD.t3127 10.4172
R2393 VDD.t4112 VDD.t205 10.4172
R2394 VDD.n1719 VDD.t3736 10.3175
R2395 VDD.n1893 VDD.t647 10.238
R2396 VDD.n145 VDD.n144 9.82175
R2397 VDD.n135 VDD.n134 9.7025
R2398 VDD.n112 VDD.t373 9.65475
R2399 VDD.t3473 VDD.t277 9.55845
R2400 VDD.t2054 VDD.t32 9.53566
R2401 VDD.t1084 VDD.t1038 9.53566
R2402 VDD.n116 VDD.t377 9.48844
R2403 VDD.n349 VDD.n342 9.45024
R2404 VDD.n2115 VDD.n2109 9.33541
R2405 VDD.t3901 VDD.t1112 9.25976
R2406 VDD.t1360 VDD.t1765 9.25976
R2407 VDD.t4148 VDD.t2109 9.25976
R2408 VDD.t3190 VDD.t2508 9.25976
R2409 VDD.t4090 VDD.t3228 9.25976
R2410 VDD.t520 VDD.t2568 9.25976
R2411 VDD.t179 VDD.t835 9.25976
R2412 VDD.t169 VDD.t839 9.25976
R2413 VDD.t167 VDD.t833 9.25976
R2414 VDD.t157 VDD.t831 9.25976
R2415 VDD.t141 VDD.t1798 9.25976
R2416 VDD.t151 VDD.t1806 9.25976
R2417 VDD.t412 VDD.t492 9.25976
R2418 VDD.n541 VDD.t1564 9.11778
R2419 VDD.n1660 VDD.t3328 9.11778
R2420 VDD.n1499 VDD.t2911 9.06272
R2421 VDD.n1485 VDD.t3561 9.06272
R2422 VDD.n1466 VDD.t3922 9.06272
R2423 VDD.n1429 VDD.t1721 9.06272
R2424 VDD.n1401 VDD.t907 9.06272
R2425 VDD.n1538 VDD.t3506 9.06272
R2426 VDD.n1567 VDD.t2982 9.06272
R2427 VDD.n1640 VDD.t3653 9.06272
R2428 VDD.n1617 VDD.t2933 9.06272
R2429 VDD.n1284 VDD.t1972 9.06272
R2430 VDD.n1289 VDD.t1780 9.06272
R2431 VDD.n1720 VDD.t2965 9.06272
R2432 VDD.n452 VDD.t2971 9.06272
R2433 VDD.n1800 VDD.t1026 9.06272
R2434 VDD.n1831 VDD.t1478 9.06272
R2435 VDD.n1105 VDD.t1198 9.06272
R2436 VDD.n1867 VDD.t1494 9.06272
R2437 VDD.n356 VDD.t3670 9.06272
R2438 VDD.n1940 VDD.t4180 9.06272
R2439 VDD.n1974 VDD.t1094 9.06272
R2440 VDD.n1998 VDD.t4031 9.06272
R2441 VDD.n2029 VDD.t2242 9.06272
R2442 VDD.n2010 VDD.t2990 9.06272
R2443 VDD.n2060 VDD.t2079 9.06272
R2444 VDD.n286 VDD.t3792 9.06272
R2445 VDD.n2047 VDD.t1978 9.06272
R2446 VDD.n2125 VDD.t938 9.06272
R2447 VDD.t2926 VDD.t513 8.80922
R2448 VDD.n117 VDD.n115 8.43844
R2449 VDD.n118 VDD.n114 8.43844
R2450 VDD.n113 VDD.n110 8.43844
R2451 VDD.n112 VDD.n111 8.43844
R2452 VDD.t769 VDD.t422 8.10235
R2453 VDD.t3324 VDD.t3931 8.10235
R2454 VDD.t2260 VDD.t912 8.10235
R2455 VDD.t2353 VDD.t876 8.10235
R2456 VDD.t2920 VDD.t3819 8.10235
R2457 VDD.n312 VDD.t411 8.0005
R2458 VDD.n1502 VDD.t3966 7.70854
R2459 VDD.n1490 VDD.t1612 7.70854
R2460 VDD.n1461 VDD.t2431 7.70854
R2461 VDD.n1434 VDD.t3880 7.70854
R2462 VDD.n1405 VDD.t2471 7.70854
R2463 VDD.n1541 VDD.t1766 7.70854
R2464 VDD.n1565 VDD.t3308 7.70854
R2465 VDD.n1636 VDD.t4029 7.70854
R2466 VDD.n1614 VDD.t3711 7.70854
R2467 VDD.n1279 VDD.t4146 7.70854
R2468 VDD.n1285 VDD.t2787 7.70854
R2469 VDD.n1725 VDD.t40 7.70854
R2470 VDD.n448 VDD.t1028 7.70854
R2471 VDD.n1797 VDD.t1526 7.70854
R2472 VDD.n1770 VDD.t1799 7.70854
R2473 VDD.n1111 VDD.t1256 7.70854
R2474 VDD.n1863 VDD.t911 7.70854
R2475 VDD.n353 VDD.t2923 7.70854
R2476 VDD.n1943 VDD.t2867 7.70854
R2477 VDD.n1970 VDD.t2177 7.70854
R2478 VDD.n1995 VDD.t2949 7.70854
R2479 VDD.n2027 VDD.t1549 7.70854
R2480 VDD.n2007 VDD.t1673 7.70854
R2481 VDD.n2064 VDD.t1414 7.70854
R2482 VDD.n282 VDD.t1534 7.70854
R2483 VDD.n2044 VDD.t2467 7.70854
R2484 VDD.n2121 VDD.t3310 7.70854
R2485 VDD.n1530 VDD.t766 7.66619
R2486 VDD.n1665 VDD.t538 7.66619
R2487 VDD.n1697 VDD.t3732 7.5363
R2488 VDD.n1713 VDD.t25 7.5363
R2489 VDD.n1727 VDD.t826 7.5061
R2490 VDD.n1765 VDD.t150 7.5061
R2491 VDD.n1771 VDD.t140 7.5061
R2492 VDD.n1823 VDD.t44 7.5061
R2493 VDD.n1822 VDD.t126 7.5061
R2494 VDD.n1179 VDD.t2000 7.5061
R2495 VDD.n1118 VDD.t444 7.5061
R2496 VDD.n2144 VDD.t2739 7.5061
R2497 VDD.n2142 VDD.t720 7.5061
R2498 VDD.n183 VDD.t332 7.50384
R2499 VDD.n178 VDD.t340 7.30419
R2500 VDD.n565 VDD.t3434 7.20842
R2501 VDD.n574 VDD.t3605 7.20842
R2502 VDD.n580 VDD.t3647 7.20842
R2503 VDD.n609 VDD.t3414 7.20842
R2504 VDD.n1397 VDD.t3282 7.20842
R2505 VDD.n523 VDD.t3348 7.20842
R2506 VDD.n501 VDD.t1829 7.20842
R2507 VDD.n1590 VDD.t3020 7.20842
R2508 VDD.n1606 VDD.t3541 7.20842
R2509 VDD.n1269 VDD.t3617 7.20842
R2510 VDD.n1266 VDD.t1154 7.20842
R2511 VDD.n421 VDD.t1528 7.20842
R2512 VDD.n442 VDD.t1862 7.20842
R2513 VDD.n1790 VDD.t2951 7.20842
R2514 VDD.n387 VDD.t3960 7.20842
R2515 VDD.n1100 VDD.t4174 7.20842
R2516 VDD.n1854 VDD.t3195 7.20842
R2517 VDD.n344 VDD.t1023 7.20842
R2518 VDD.n315 VDD.t1520 7.20842
R2519 VDD.n1959 VDD.t995 7.20842
R2520 VDD.n1942 VDD.t4008 7.20842
R2521 VDD.n292 VDD.t3691 7.20842
R2522 VDD.n300 VDD.t2060 7.20842
R2523 VDD.n259 VDD.t1625 7.20842
R2524 VDD.n271 VDD.t1570 7.20842
R2525 VDD.n261 VDD.t2684 7.20842
R2526 VDD.n2108 VDD.t2828 7.20842
R2527 VDD.n537 VDD.t6 7.18658
R2528 VDD.n1625 VDD.t797 7.18658
R2529 VDD.n479 VDD.t3225 7.18658
R2530 VDD.n450 VDD.t4142 7.18658
R2531 VDD.n354 VDD.t1096 7.18658
R2532 VDD.n1939 VDD.t3090 7.18658
R2533 VDD.n2026 VDD.t4206 7.18658
R2534 VDD.n2039 VDD.t2969 7.18658
R2535 VDD.n2134 VDD.t3274 7.18658
R2536 VDD.n527 VDD.t1897 7.17999
R2537 VDD.n467 VDD.t4231 7.17999
R2538 VDD.t2981 VDD.n502 7.16896
R2539 VDD.n1419 VDD.n636 7.15066
R2540 VDD.n680 VDD.n214 7.15066
R2541 VDD.n2333 VDD.n215 7.15066
R2542 VDD.n1524 VDD.n546 7.15066
R2543 VDD.n535 VDD.t438 7.01851
R2544 VDD.n1627 VDD.t3430 7.01851
R2545 VDD.n1646 VDD.t2905 7.01851
R2546 VDD.n449 VDD.t2519 7.01851
R2547 VDD.n351 VDD.t2741 7.01851
R2548 VDD.n1938 VDD.t2848 7.01851
R2549 VDD.n2024 VDD.t3639 7.01851
R2550 VDD.n2041 VDD.t3276 7.01851
R2551 VDD.n2135 VDD.t3589 7.01851
R2552 VDD.n562 VDD.t891 7.0005
R2553 VDD.n1374 VDD.t2651 7.0005
R2554 VDD.n1388 VDD.t2110 7.0005
R2555 VDD.n507 VDD.t3448 7.0005
R2556 VDD.n508 VDD.t3055 7.0005
R2557 VDD.n513 VDD.t3261 7.0005
R2558 VDD.n1387 VDD.t1271 7.0005
R2559 VDD.n1343 VDD.t1710 7.0005
R2560 VDD.n1349 VDD.t2132 7.0005
R2561 VDD.n489 VDD.t1348 7.0005
R2562 VDD.n1602 VDD.t3191 7.0005
R2563 VDD.n1605 VDD.t4223 7.0005
R2564 VDD.n1603 VDD.t1926 7.0005
R2565 VDD.n1599 VDD.t3781 7.0005
R2566 VDD.n488 VDD.t1955 7.0005
R2567 VDD.n1263 VDD.t2762 7.0005
R2568 VDD.n466 VDD.t3483 7.0005
R2569 VDD.n440 VDD.t1335 7.0005
R2570 VDD.n439 VDD.t3762 7.0005
R2571 VDD.n1176 VDD.t1145 7.0005
R2572 VDD.n1789 VDD.t2567 7.0005
R2573 VDD.n369 VDD.t1115 7.0005
R2574 VDD.n372 VDD.t2881 7.0005
R2575 VDD.n1099 VDD.t1555 7.0005
R2576 VDD.n327 VDD.t2146 7.0005
R2577 VDD.n337 VDD.t956 7.0005
R2578 VDD.n343 VDD.t3855 7.0005
R2579 VDD.n340 VDD.t2235 7.0005
R2580 VDD.n326 VDD.t2656 7.0005
R2581 VDD.n1952 VDD.t1736 7.0005
R2582 VDD.n1955 VDD.t1949 7.0005
R2583 VDD.n921 VDD.t3704 7.0005
R2584 VDD.n299 VDD.t3176 7.0005
R2585 VDD.n2019 VDD.t2589 7.0005
R2586 VDD.n920 VDD.t879 7.0005
R2587 VDD.n268 VDD.t1185 7.0005
R2588 VDD.n256 VDD.t1579 7.0005
R2589 VDD.n2106 VDD.t3502 7.0005
R2590 VDD.n1280 VDD.t1045 6.88796
R2591 VDD.n1591 VDD.t2053 6.88404
R2592 VDD.n1688 VDD.t1893 6.88404
R2593 VDD.n304 VDD.t237 6.8755
R2594 VDD.n1637 VDD.t3510 6.84883
R2595 VDD.n1581 VDD.t2806 6.84883
R2596 VDD.n2137 VDD.t4196 6.84883
R2597 VDD.n1554 VDD.t1391 6.80877
R2598 VDD.n1587 VDD.t1273 6.80877
R2599 VDD.n1657 VDD.t3257 6.80877
R2600 VDD.n1897 VDD.t3676 6.80877
R2601 VDD.n1902 VDD.t1053 6.80877
R2602 VDD.n527 VDD.t2909 6.31276
R2603 VDD.n467 VDD.t3633 6.31276
R2604 VDD.n183 VDD.n182 6.25419
R2605 VDD.n184 VDD.n181 6.25419
R2606 VDD.n180 VDD.n176 6.25419
R2607 VDD.n179 VDD.n177 6.25419
R2608 VDD.t2983 VDD.t794 5.97422
R2609 VDD.n575 VDD.t4025 5.9474
R2610 VDD.n547 VDD.t2185 5.9474
R2611 VDD.n496 VDD.t1032 5.9474
R2612 VDD.n1348 VDD.t138 5.9474
R2613 VDD.n1347 VDD.t3463 5.9474
R2614 VDD.n360 VDD.t845 5.9474
R2615 VDD.n317 VDD.t4153 5.9474
R2616 VDD.n313 VDD.t3984 5.9474
R2617 VDD.n917 VDD.t2314 5.9474
R2618 VDD.n2110 VDD.t1324 5.9474
R2619 VDD.n1286 VDD.n1269 5.90374
R2620 VDD.n1716 VDD.n421 5.90374
R2621 VDD.n1498 VDD.n565 5.89642
R2622 VDD.n1480 VDD.n574 5.89642
R2623 VDD.n1469 VDD.n580 5.89642
R2624 VDD.n1426 VDD.n609 5.89642
R2625 VDD.n1399 VDD.n1397 5.89642
R2626 VDD.n1534 VDD.n523 5.89642
R2627 VDD.n1571 VDD.n501 5.89642
R2628 VDD.n1592 VDD.n1590 5.89642
R2629 VDD.n1619 VDD.n1606 5.89642
R2630 VDD.n1293 VDD.n1266 5.89642
R2631 VDD.n455 VDD.n442 5.89642
R2632 VDD.n1802 VDD.n1790 5.89642
R2633 VDD.n1828 VDD.n387 5.89642
R2634 VDD.n1102 VDD.n1100 5.89642
R2635 VDD.n1855 VDD.n1854 5.89642
R2636 VDD.n358 VDD.n344 5.89642
R2637 VDD.n1937 VDD.n315 5.89642
R2638 VDD.n1978 VDD.n1959 5.89642
R2639 VDD.n1944 VDD.n1942 5.89642
R2640 VDD.n293 VDD.n292 5.89642
R2641 VDD.n2012 VDD.n300 5.89642
R2642 VDD.n2057 VDD.n259 5.89642
R2643 VDD.n290 VDD.n271 5.89642
R2644 VDD.n2051 VDD.n261 5.89642
R2645 VDD.n2128 VDD.n2108 5.89642
R2646 VDD.n425 VDD.t1043 5.79932
R2647 VDD.n422 VDD.t1041 5.79932
R2648 VDD.t3083 VDD.t3504 5.78754
R2649 VDD.t2766 VDD.t3400 5.78754
R2650 VDD.t2987 VDD.n1386 5.78754
R2651 VDD.t2761 VDD.t1160 5.78754
R2652 VDD.t2647 VDD.t1144 5.78754
R2653 VDD.t3677 VDD.t3955 5.78754
R2654 VDD.t485 VDD.t1773 5.78754
R2655 VDD.t530 VDD.t1622 5.78754
R2656 VDD.n1533 VDD.n524 5.55267
R2657 VDD.n458 VDD.n457 5.55267
R2658 VDD.n350 VDD.n348 5.45352
R2659 VDD.n563 VDD.t722 5.38512
R2660 VDD.n571 VDD.t709 5.38512
R2661 VDD.n584 VDD.t755 5.38512
R2662 VDD.n606 VDD.t764 5.38512
R2663 VDD.n1394 VDD.t714 5.38512
R2664 VDD.n521 VDD.t757 5.38512
R2665 VDD.n503 VDD.t748 5.38512
R2666 VDD.n484 VDD.t532 5.38512
R2667 VDD.n1608 VDD.t468 5.38512
R2668 VDD.n1271 VDD.t774 5.38512
R2669 VDD.n1268 VDD.t750 5.38512
R2670 VDD.n418 VDD.t702 5.38512
R2671 VDD.n444 VDD.t528 5.38512
R2672 VDD.n1793 VDD.t476 5.38512
R2673 VDD.n383 VDD.t482 5.38512
R2674 VDD.n1096 VDD.t752 5.38512
R2675 VDD.n364 VDD.t478 5.38512
R2676 VDD.n346 VDD.t474 5.38512
R2677 VDD.n1941 VDD.t724 5.38512
R2678 VDD.n1963 VDD.t518 5.38512
R2679 VDD.n311 VDD.t493 5.38512
R2680 VDD.n295 VDD.t462 5.38512
R2681 VDD.n302 VDD.t484 5.38512
R2682 VDD.n257 VDD.t535 5.38512
R2683 VDD.n275 VDD.t498 5.38512
R2684 VDD.n264 VDD.t491 5.38512
R2685 VDD.n2111 VDD.t508 5.38512
R2686 VDD.n1652 VDD.n474 5.38246
R2687 VDD.n1649 VDD.n475 5.38246
R2688 VDD.n1647 VDD.n477 5.38246
R2689 VDD.n1645 VDD.n478 5.38246
R2690 VDD.n1275 VDD.n1274 5.38246
R2691 VDD.n1698 VDD.n433 5.38246
R2692 VDD.n1700 VDD.n431 5.38246
R2693 VDD.n1702 VDD.n429 5.38246
R2694 VDD.n1704 VDD.n427 5.38246
R2695 VDD.n1706 VDD.n425 5.38246
R2696 VDD.n1708 VDD.n423 5.38246
R2697 VDD.n1711 VDD.n422 5.38246
R2698 VDD.n1504 VDD.n561 5.36991
R2699 VDD.n1492 VDD.n567 5.36991
R2700 VDD.n1459 VDD.n587 5.36991
R2701 VDD.n1436 VDD.n602 5.36991
R2702 VDD.n1407 VDD.n1392 5.36991
R2703 VDD.n1543 VDD.n518 5.36991
R2704 VDD.n1563 VDD.n505 5.36991
R2705 VDD.n1634 VDD.n486 5.36991
R2706 VDD.n1612 VDD.n1611 5.36991
R2707 VDD.n1276 VDD.n1273 5.36991
R2708 VDD.n1283 VDD.n1270 5.36991
R2709 VDD.n1728 VDD.n416 5.36991
R2710 VDD.n447 VDD.n445 5.36991
R2711 VDD.n1796 VDD.n1794 5.36991
R2712 VDD.n1772 VDD.n1769 5.36991
R2713 VDD.n1113 VDD.n1092 5.36991
R2714 VDD.n1861 VDD.n367 5.36991
R2715 VDD.n352 VDD.n347 5.36991
R2716 VDD.n310 VDD.n309 5.36991
R2717 VDD.n1968 VDD.n1966 5.36991
R2718 VDD.n1993 VDD.n314 5.36991
R2719 VDD.n2025 VDD.n296 5.36991
R2720 VDD.n2005 VDD.n305 5.36991
R2721 VDD.n2066 VDD.n254 5.36991
R2722 VDD.n280 VDD.n278 5.36991
R2723 VDD.n2042 VDD.n267 5.36991
R2724 VDD.n2119 VDD.n2113 5.36991
R2725 VDD.n627 VDD.n617 5.36093
R2726 VDD.n629 VDD.n615 5.36093
R2727 VDD.n631 VDD.n613 5.36093
R2728 VDD.n1421 VDD.n611 5.36093
R2729 VDD.n1428 VDD.n608 5.36093
R2730 VDD.n1430 VDD.n607 5.36093
R2731 VDD.n1432 VDD.n605 5.36093
R2732 VDD.n1435 VDD.n603 5.36093
R2733 VDD.n1448 VDD.n595 5.36093
R2734 VDD.n1450 VDD.n593 5.36093
R2735 VDD.n1453 VDD.n591 5.36093
R2736 VDD.n1457 VDD.n588 5.36093
R2737 VDD.n1465 VDD.n583 5.36093
R2738 VDD.n1467 VDD.n582 5.36093
R2739 VDD.n1468 VDD.n581 5.36093
R2740 VDD.n1473 VDD.n578 5.36093
R2741 VDD.n1484 VDD.n573 5.36093
R2742 VDD.n1486 VDD.n572 5.36093
R2743 VDD.n1488 VDD.n570 5.36093
R2744 VDD.n1491 VDD.n568 5.36093
R2745 VDD.n1522 VDD.n549 5.36093
R2746 VDD.n1518 VDD.n552 5.36093
R2747 VDD.n1516 VDD.n554 5.36093
R2748 VDD.n1514 VDD.n556 5.36093
R2749 VDD.n1511 VDD.n558 5.36093
R2750 VDD.n1513 VDD.n557 5.36093
R2751 VDD.n1515 VDD.n555 5.36093
R2752 VDD.n1519 VDD.n551 5.36093
R2753 VDD.n1451 VDD.n592 5.36093
R2754 VDD.n1447 VDD.n596 5.36093
R2755 VDD.n1445 VDD.n597 5.36093
R2756 VDD.n1443 VDD.n599 5.36093
R2757 VDD.n630 VDD.n614 5.36093
R2758 VDD.n626 VDD.n618 5.36093
R2759 VDD.n624 VDD.n619 5.36093
R2760 VDD.n622 VDD.n620 5.36093
R2761 VDD.n536 VDD.n533 5.36093
R2762 VDD.n538 VDD.n532 5.36093
R2763 VDD.n540 VDD.n530 5.36093
R2764 VDD.n543 VDD.n528 5.36093
R2765 VDD.n1677 VDD.n460 5.36093
R2766 VDD.n1672 VDD.n464 5.36093
R2767 VDD.n1674 VDD.n463 5.36093
R2768 VDD.n1675 VDD.n462 5.36093
R2769 VDD.n1678 VDD.n459 5.36093
R2770 VDD.n1655 VDD.n472 5.36093
R2771 VDD.n1696 VDD.n434 5.36093
R2772 VDD.n453 VDD.n443 5.36093
R2773 VDD.n1860 VDD.n368 5.36093
R2774 VDD.n1862 VDD.n366 5.36093
R2775 VDD.n1864 VDD.n365 5.36093
R2776 VDD.n1868 VDD.n362 5.36093
R2777 VDD.n1884 VDD.n335 5.36093
R2778 VDD.n1990 VDD.n1951 5.36093
R2779 VDD.n1969 VDD.n1965 5.36093
R2780 VDD.n1971 VDD.n1964 5.36093
R2781 VDD.n1973 VDD.n1962 5.36093
R2782 VDD.n1976 VDD.n1960 5.36093
R2783 VDD.n1985 VDD.n1956 5.36093
R2784 VDD.n2003 VDD.n306 5.36093
R2785 VDD.n2016 VDD.n298 5.36093
R2786 VDD.n2054 VDD.n260 5.36093
R2787 VDD.n281 VDD.n277 5.36093
R2788 VDD.n283 VDD.n276 5.36093
R2789 VDD.n285 VDD.n274 5.36093
R2790 VDD.n288 VDD.n272 5.36093
R2791 VDD.n2177 VDD.n236 5.36093
R2792 VDD.n2179 VDD.n235 5.36093
R2793 VDD.n2181 VDD.n234 5.36093
R2794 VDD.n2185 VDD.n232 5.36093
R2795 VDD.n2289 VDD.n2286 5.36093
R2796 VDD.n2291 VDD.n2285 5.36093
R2797 VDD.n2293 VDD.n2284 5.36093
R2798 VDD.n2297 VDD.n2282 5.36093
R2799 VDD.n1729 VDD.n415 5.35702
R2800 VDD.n1732 VDD.n412 5.35702
R2801 VDD.n1734 VDD.n410 5.35702
R2802 VDD.n1736 VDD.n408 5.35702
R2803 VDD.n1755 VDD.n397 5.35702
R2804 VDD.n1757 VDD.n395 5.35702
R2805 VDD.n1759 VDD.n393 5.35702
R2806 VDD.n1763 VDD.n389 5.35702
R2807 VDD.n381 VDD.n380 5.35702
R2808 VDD.n1832 VDD.n384 5.35702
R2809 VDD.n1830 VDD.n385 5.35702
R2810 VDD.n1829 VDD.n386 5.35702
R2811 VDD.n1821 VDD.n1777 5.35702
R2812 VDD.n1817 VDD.n1781 5.35702
R2813 VDD.n1815 VDD.n1783 5.35702
R2814 VDD.n1813 VDD.n1785 5.35702
R2815 VDD.n1812 VDD.n1786 5.35702
R2816 VDD.n1814 VDD.n1784 5.35702
R2817 VDD.n1816 VDD.n1782 5.35702
R2818 VDD.n1820 VDD.n1778 5.35702
R2819 VDD.n1747 VDD.n402 5.35702
R2820 VDD.n1745 VDD.n403 5.35702
R2821 VDD.n405 VDD.n404 5.35702
R2822 VDD.n1109 VDD.n1095 5.35702
R2823 VDD.n1110 VDD.n1094 5.35702
R2824 VDD.n1112 VDD.n1093 5.35702
R2825 VDD.n1117 VDD.n1090 5.35702
R2826 VDD.n2100 VDD.n2099 5.35702
R2827 VDD.n243 VDD.n241 5.35702
R2828 VDD.n243 VDD.n242 5.35702
R2829 VDD.n2148 VDD.n244 5.35702
R2830 VDD.n2148 VDD.n245 5.35702
R2831 VDD.n2147 VDD.n247 5.35702
R2832 VDD.n2145 VDD.n249 5.35702
R2833 VDD.n2144 VDD.n250 5.35702
R2834 VDD.n539 VDD.n531 5.35271
R2835 VDD.n1658 VDD.n470 5.35271
R2836 VDD.n1546 VDD.n516 5.34344
R2837 VDD.n1540 VDD.n520 5.34344
R2838 VDD.n1558 VDD.n509 5.34344
R2839 VDD.n1400 VDD.n1396 5.34344
R2840 VDD.n1360 VDD.n1344 5.34344
R2841 VDD.n1773 VDD.n1768 5.34344
R2842 VDD.n1844 VDD.n374 5.34344
R2843 VDD.n1501 VDD.n563 5.33285
R2844 VDD.n1487 VDD.n571 5.33285
R2845 VDD.n1464 VDD.n584 5.33285
R2846 VDD.n1431 VDD.n606 5.33285
R2847 VDD.n1403 VDD.n1394 5.33285
R2848 VDD.n1539 VDD.n521 5.33285
R2849 VDD.n1566 VDD.n503 5.33285
R2850 VDD.n1638 VDD.n484 5.33285
R2851 VDD.n1616 VDD.n1608 5.33285
R2852 VDD.n1282 VDD.n1271 5.33285
R2853 VDD.n1287 VDD.n1268 5.33285
R2854 VDD.n1722 VDD.n418 5.33285
R2855 VDD.n451 VDD.n444 5.33285
R2856 VDD.n1798 VDD.n1793 5.33285
R2857 VDD.n1833 VDD.n383 5.33285
R2858 VDD.n1108 VDD.n1096 5.33285
R2859 VDD.n1865 VDD.n364 5.33285
R2860 VDD.n355 VDD.n346 5.33285
R2861 VDD.n1947 VDD.n1941 5.33285
R2862 VDD.n1972 VDD.n1963 5.33285
R2863 VDD.n1997 VDD.n311 5.33285
R2864 VDD.n2028 VDD.n295 5.33285
R2865 VDD.n2009 VDD.n302 5.33285
R2866 VDD.n2061 VDD.n257 5.33285
R2867 VDD.n284 VDD.n275 5.33285
R2868 VDD.n2046 VDD.n264 5.33285
R2869 VDD.n2123 VDD.n2111 5.33285
R2870 VDD.n1707 VDD.n424 5.31789
R2871 VDD.n1555 VDD.n512 5.31697
R2872 VDD.n1589 VDD.n487 5.31697
R2873 VDD.n1656 VDD.n471 5.31697
R2874 VDD.n1894 VDD.n329 5.31697
R2875 VDD.n1903 VDD.n323 5.31697
R2876 VDD.n1639 VDD.n483 5.30638
R2877 VDD.n1579 VDD.n495 5.30638
R2878 VDD.n2139 VDD.n2105 5.30638
R2879 VDD.n1721 VDD.n419 5.30615
R2880 VDD.n1723 VDD.n417 5.30615
R2881 VDD.n1891 VDD.n331 5.30615
R2882 VDD.n1889 VDD.n333 5.30615
R2883 VDD.n1537 VDD.n522 5.29976
R2884 VDD.n1648 VDD.n476 5.29976
R2885 VDD.n1667 VDD.n1666 5.29976
R2886 VDD.n2048 VDD.n263 5.29976
R2887 VDD.n1444 VDD.n598 5.28785
R2888 VDD.n1462 VDD.n585 5.28785
R2889 VDD.n1500 VDD.n564 5.28785
R2890 VDD.n1510 VDD.n559 5.28785
R2891 VDD.n1456 VDD.n589 5.28785
R2892 VDD.n1380 VDD.n1375 5.28785
R2893 VDD.n1410 VDD.n1390 5.28785
R2894 VDD.n1564 VDD.n504 5.28785
R2895 VDD.n1556 VDD.n511 5.28785
R2896 VDD.n1528 VDD.n526 5.28785
R2897 VDD.n1547 VDD.n515 5.28785
R2898 VDD.n1408 VDD.n1391 5.28785
R2899 VDD.n1412 VDD.n1389 5.28785
R2900 VDD.n1366 VDD.n1341 5.28785
R2901 VDD.n1358 VDD.n1345 5.28785
R2902 VDD.n1352 VDD.n1351 5.28785
R2903 VDD.n1583 VDD.n492 5.28785
R2904 VDD.n1630 VDD.n1600 5.28785
R2905 VDD.n1613 VDD.n1610 5.28785
R2906 VDD.n1615 VDD.n1609 5.28785
R2907 VDD.n1629 VDD.n1601 5.28785
R2908 VDD.n1635 VDD.n485 5.28785
R2909 VDD.n482 VDD.n481 5.28785
R2910 VDD.n1585 VDD.n490 5.28785
R2911 VDD.n1584 VDD.n491 5.28785
R2912 VDD.n1582 VDD.n493 5.28785
R2913 VDD.n498 VDD.n497 5.28785
R2914 VDD.n1353 VDD.n1350 5.28785
R2915 VDD.n1304 VDD.n1264 5.28785
R2916 VDD.n1671 VDD.n465 5.28785
R2917 VDD.n1661 VDD.n468 5.28785
R2918 VDD.n1659 VDD.n469 5.28785
R2919 VDD.n1733 VDD.n411 5.28785
R2920 VDD.n1730 VDD.n414 5.28785
R2921 VDD.n1694 VDD.n436 5.28785
R2922 VDD.n1692 VDD.n438 5.28785
R2923 VDD.n447 VDD.n446 5.28785
R2924 VDD.n1695 VDD.n435 5.28785
R2925 VDD.n1178 VDD.n1177 5.28785
R2926 VDD.n1799 VDD.n1792 5.28785
R2927 VDD.n1801 VDD.n1791 5.28785
R2928 VDD.n1808 VDD.n1787 5.28785
R2929 VDD.n1849 VDD.n371 5.28785
R2930 VDD.n1850 VDD.n370 5.28785
R2931 VDD.n1842 VDD.n375 5.28785
R2932 VDD.n1839 VDD.n377 5.28785
R2933 VDD.n1904 VDD.n322 5.28785
R2934 VDD.n1901 VDD.n324 5.28785
R2935 VDD.n1880 VDD.n339 5.28785
R2936 VDD.n1878 VDD.n341 5.28785
R2937 VDD.n357 VDD.n345 5.28785
R2938 VDD.n1883 VDD.n336 5.28785
R2939 VDD.n1890 VDD.n332 5.28785
R2940 VDD.n1892 VDD.n330 5.28785
R2941 VDD.n1895 VDD.n328 5.28785
R2942 VDD.n1905 VDD.n321 5.28785
R2943 VDD.n1987 VDD.n1954 5.28785
R2944 VDD.n1981 VDD.n1958 5.28785
R2945 VDD.n1988 VDD.n1953 5.28785
R2946 VDD.n1933 VDD.n316 5.28785
R2947 VDD.n929 VDD.n916 5.28785
R2948 VDD.n2011 VDD.n301 5.28785
R2949 VDD.n2017 VDD.n297 5.28785
R2950 VDD.n2030 VDD.n294 5.28785
R2951 VDD.n923 VDD.n922 5.28785
R2952 VDD.n2045 VDD.n265 5.28785
R2953 VDD.n2035 VDD.n270 5.28785
R2954 VDD.n2059 VDD.n258 5.28785
R2955 VDD.n2122 VDD.n2112 5.28785
R2956 VDD.n2132 VDD.n2107 5.28785
R2957 VDD.n2171 VDD.n237 5.28785
R2958 VDD.n2315 VDD.n2280 5.28785
R2959 VDD.n1731 VDD.n413 5.28659
R2960 VDD.n1761 VDD.n391 5.28659
R2961 VDD.n1834 VDD.n382 5.28659
R2962 VDD.n1819 VDD.n1779 5.28659
R2963 VDD.n1818 VDD.n1780 5.28659
R2964 VDD.n1764 VDD.n388 5.28659
R2965 VDD.n1762 VDD.n390 5.28659
R2966 VDD.n1760 VDD.n392 5.28659
R2967 VDD.n1758 VDD.n394 5.28659
R2968 VDD.n1756 VDD.n396 5.28659
R2969 VDD.n1754 VDD.n398 5.28659
R2970 VDD.n1751 VDD.n399 5.28659
R2971 VDD.n1749 VDD.n400 5.28659
R2972 VDD.n1115 VDD.n1091 5.28659
R2973 VDD.n2147 VDD.n246 5.28659
R2974 VDD.n2146 VDD.n248 5.28659
R2975 VDD.n1479 VDD.n575 5.27991
R2976 VDD.n548 VDD.n547 5.27991
R2977 VDD.n1578 VDD.n496 5.27991
R2978 VDD.n1355 VDD.n1348 5.27991
R2979 VDD.n1356 VDD.n1347 5.27991
R2980 VDD.n361 VDD.n360 5.27991
R2981 VDD.n1932 VDD.n317 5.27991
R2982 VDD.n1994 VDD.n313 5.27991
R2983 VDD.n928 VDD.n917 5.27991
R2984 VDD.n2126 VDD.n2110 5.27991
R2985 VDD.n1503 VDD.n562 5.25874
R2986 VDD.n1383 VDD.n1374 5.25874
R2987 VDD.n1413 VDD.n1388 5.25874
R2988 VDD.n1560 VDD.n507 5.25874
R2989 VDD.n1559 VDD.n508 5.25874
R2990 VDD.n1552 VDD.n513 5.25874
R2991 VDD.n1415 VDD.n1387 5.25874
R2992 VDD.n1361 VDD.n1343 5.25874
R2993 VDD.n1354 VDD.n1349 5.25874
R2994 VDD.n1586 VDD.n489 5.25874
R2995 VDD.n1628 VDD.n1602 5.25874
R2996 VDD.n1618 VDD.n1607 5.25874
R2997 VDD.n1621 VDD.n1605 5.25874
R2998 VDD.n1626 VDD.n1603 5.25874
R2999 VDD.n1632 VDD.n1599 5.25874
R3000 VDD.n1588 VDD.n488 5.25874
R3001 VDD.n1305 VDD.n1263 5.25874
R3002 VDD.n1664 VDD.n466 5.25874
R3003 VDD.n1705 VDD.n426 5.25874
R3004 VDD.n1703 VDD.n428 5.25874
R3005 VDD.n1701 VDD.n430 5.25874
R3006 VDD.n1690 VDD.n440 5.25874
R3007 VDD.n1691 VDD.n439 5.25874
R3008 VDD.n1693 VDD.n437 5.25874
R3009 VDD.n1180 VDD.n1176 5.25874
R3010 VDD.n1804 VDD.n1789 5.25874
R3011 VDD.n1851 VDD.n369 5.25874
R3012 VDD.n1848 VDD.n372 5.25874
R3013 VDD.n1103 VDD.n1099 5.25874
R3014 VDD.n1898 VDD.n327 5.25874
R3015 VDD.n1882 VDD.n337 5.25874
R3016 VDD.n1874 VDD.n343 5.25874
R3017 VDD.n1879 VDD.n340 5.25874
R3018 VDD.n1881 VDD.n338 5.25874
R3019 VDD.n1899 VDD.n326 5.25874
R3020 VDD.n1989 VDD.n1952 5.25874
R3021 VDD.n1986 VDD.n1955 5.25874
R3022 VDD.n927 VDD.n918 5.25874
R3023 VDD.n924 VDD.n921 5.25874
R3024 VDD.n2015 VDD.n299 5.25874
R3025 VDD.n2020 VDD.n2019 5.25874
R3026 VDD.n925 VDD.n920 5.25874
R3027 VDD.n2043 VDD.n266 5.25874
R3028 VDD.n2040 VDD.n268 5.25874
R3029 VDD.n2062 VDD.n256 5.25874
R3030 VDD.n2136 VDD.n2106 5.25874
R3031 VDD.n524 VDD.t3139 5.20563
R3032 VDD.n457 VDD.t2688 5.20563
R3033 VDD.n1846 VDD.t3581 5.15426
R3034 VDD.n1887 VDD.t1917 5.15426
R3035 VDD.n564 VDD.t2075 5.05606
R3036 VDD.n562 VDD.t1706 5.05606
R3037 VDD.n1374 VDD.t2767 5.05606
R3038 VDD.n1375 VDD.t2732 5.05606
R3039 VDD.n1388 VDD.t2169 5.05606
R3040 VDD.n1390 VDD.t1849 5.05606
R3041 VDD.n504 VDD.t2105 5.05606
R3042 VDD.n507 VDD.t1545 5.05606
R3043 VDD.n508 VDD.t2187 5.05606
R3044 VDD.n511 VDD.t4252 5.05606
R3045 VDD.n515 VDD.t3323 5.05606
R3046 VDD.n513 VDD.t1447 5.05606
R3047 VDD.n1389 VDD.t4149 5.05606
R3048 VDD.n1387 VDD.t2988 5.05606
R3049 VDD.n1343 VDD.t2973 5.05606
R3050 VDD.n1345 VDD.t3548 5.05606
R3051 VDD.n1349 VDD.t1604 5.05606
R3052 VDD.n1351 VDD.t1952 5.05606
R3053 VDD.n492 VDD.t1397 5.05606
R3054 VDD.n489 VDD.t2542 5.05606
R3055 VDD.n1600 VDD.t3115 5.05606
R3056 VDD.n1602 VDD.t156 5.05606
R3057 VDD.n1609 VDD.t4037 5.05606
R3058 VDD.n1607 VDD.t2200 5.05606
R3059 VDD.n1605 VDD.t2931 5.05606
R3060 VDD.n1603 VDD.t2409 5.05606
R3061 VDD.n1601 VDD.t2509 5.05606
R3062 VDD.n1599 VDD.t3767 5.05606
R3063 VDD.n485 VDD.t1484 5.05606
R3064 VDD.n488 VDD.t606 5.05606
R3065 VDD.n490 VDD.t3445 5.05606
R3066 VDD.n1263 VDD.t3461 5.05606
R3067 VDD.n1264 VDD.t2749 5.05606
R3068 VDD.n466 VDD.t1165 5.05606
R3069 VDD.n468 VDD.t1615 5.05606
R3070 VDD.n438 VDD.t2594 5.05606
R3071 VDD.n440 VDD.t2247 5.05606
R3072 VDD.n439 VDD.t3759 5.05606
R3073 VDD.n437 VDD.t1886 5.05606
R3074 VDD.n435 VDD.t1156 5.05606
R3075 VDD.n1176 VDD.t847 5.05606
R3076 VDD.n1177 VDD.t2164 5.05606
R3077 VDD.n1791 VDD.t922 5.05606
R3078 VDD.n1789 VDD.t2020 5.05606
R3079 VDD.n371 VDD.t2453 5.05606
R3080 VDD.n369 VDD.t4047 5.05606
R3081 VDD.n370 VDD.t981 5.05606
R3082 VDD.n372 VDD.t1327 5.05606
R3083 VDD.n377 VDD.t3974 5.05606
R3084 VDD.n1099 VDD.t2529 5.05606
R3085 VDD.n324 VDD.t3518 5.05606
R3086 VDD.n327 VDD.t2041 5.05606
R3087 VDD.n337 VDD.t2111 5.05606
R3088 VDD.n339 VDD.t2927 5.05606
R3089 VDD.n345 VDD.t1932 5.05606
R3090 VDD.n343 VDD.t1981 5.05606
R3091 VDD.n340 VDD.t997 5.05606
R3092 VDD.n338 VDD.t3459 5.05606
R3093 VDD.n336 VDD.t3289 5.05606
R3094 VDD.n328 VDD.t2213 5.05606
R3095 VDD.n326 VDD.t2842 5.05606
R3096 VDD.n1952 VDD.t2098 5.05606
R3097 VDD.n1954 VDD.t1542 5.05606
R3098 VDD.n1955 VDD.t1404 5.05606
R3099 VDD.n1953 VDD.t3571 5.05606
R3100 VDD.n916 VDD.t3078 5.05606
R3101 VDD.n918 VDD.t3185 5.05606
R3102 VDD.n921 VDD.t2089 5.05606
R3103 VDD.n301 VDD.t2855 5.05606
R3104 VDD.n299 VDD.t4241 5.05606
R3105 VDD.n294 VDD.t1194 5.05606
R3106 VDD.n2019 VDD.t1868 5.05606
R3107 VDD.n922 VDD.t4298 5.05606
R3108 VDD.n920 VDD.t2310 5.05606
R3109 VDD.n265 VDD.t2460 5.05606
R3110 VDD.n266 VDD.t4259 5.05606
R3111 VDD.n268 VDD.t1141 5.05606
R3112 VDD.n258 VDD.t2479 5.05606
R3113 VDD.n256 VDD.t3128 5.05606
R3114 VDD.n2107 VDD.t1882 5.05606
R3115 VDD.n2106 VDD.t2429 5.05606
R3116 VDD.n1595 VDD.t3512 4.89499
R3117 VDD.n454 VDD.t1065 4.89499
R3118 VDD.n1536 VDD.t1073 4.70061
R3119 VDD.n1650 VDD.t781 4.70061
R3120 VDD.n1681 VDD.t3223 4.70061
R3121 VDD.n2049 VDD.t2259 4.70061
R3122 VDD.n1496 VDD.t3376 4.66507
R3123 VDD.n1478 VDD.t1254 4.66507
R3124 VDD.n1471 VDD.t1001 4.66507
R3125 VDD.n1423 VDD.t1574 4.66507
R3126 VDD.n1573 VDD.t1182 4.66507
R3127 VDD.n1532 VDD.t1353 4.66507
R3128 VDD.n500 VDD.t1713 4.66507
R3129 VDD.n1593 VDD.t2354 4.66507
R3130 VDD.n1622 VDD.t1974 4.66507
R3131 VDD.n1295 VDD.t1553 4.66507
R3132 VDD.n1686 VDD.t2016 4.66507
R3133 VDD.n1805 VDD.t3040 4.66507
R3134 VDD.n1826 VDD.t2907 4.66507
R3135 VDD.n1101 VDD.t1551 4.66507
R3136 VDD.n1853 VDD.t2383 4.66507
R3137 VDD.n1875 VDD.t1678 4.66507
R3138 VDD.n1936 VDD.t3467 4.66507
R3139 VDD.n1980 VDD.t1936 4.66507
R3140 VDD.n1945 VDD.t3048 4.66507
R3141 VDD.n2021 VDD.t2925 4.66507
R3142 VDD.n2013 VDD.t3888 4.66507
R3143 VDD.n2056 VDD.t2504 4.66507
R3144 VDD.n2036 VDD.t4217 4.66507
R3145 VDD.n2052 VDD.t2565 4.66507
R3146 VDD.n2129 VDD.t1909 4.66507
R3147 VDD.n1724 VDD.t1080 4.65756
R3148 VDD.n1888 VDD.t652 4.65756
R3149 VDD.t691 VDD.t864 4.63013
R3150 VDD.t3073 VDD.t920 4.63013
R3151 VDD.t85 VDD.t4045 4.63013
R3152 VDD.t307 VDD.t1879 4.63013
R3153 VDD.t1918 VDD.t3848 4.63013
R3154 VDD.n1653 VDD.t803 4.62626
R3155 VDD.n1277 VDD.t614 4.62626
R3156 VDD.t955 VDD.t2926 4.61459
R3157 VDD.n400 VDD.t1817 4.61026
R3158 VDD.n1420 VDD.n1419 4.5005
R3159 VDD.n1418 VDD.n1417 4.5005
R3160 VDD.n1372 VDD.n1371 4.5005
R3161 VDD.n1332 VDD.n1331 4.5005
R3162 VDD.n1247 VDD.n1246 4.5005
R3163 VDD.n1206 VDD.n1205 4.5005
R3164 VDD.n1160 VDD.n1159 4.5005
R3165 VDD.n1074 VDD.n1073 4.5005
R3166 VDD.n1027 VDD.n1026 4.5005
R3167 VDD.n980 VDD.n979 4.5005
R3168 VDD.n900 VDD.n899 4.5005
R3169 VDD.n853 VDD.n852 4.5005
R3170 VDD.n806 VDD.n805 4.5005
R3171 VDD.n727 VDD.n726 4.5005
R3172 VDD.n2191 VDD.n2190 4.5005
R3173 VDD.n2189 VDD.n2188 4.5005
R3174 VDD.n2124 VDD.n230 4.5005
R3175 VDD.n2034 VDD.n2033 4.5005
R3176 VDD.n2032 VDD.n2031 4.5005
R3177 VDD.n1979 VDD.n291 4.5005
R3178 VDD.n1873 VDD.n1872 4.5005
R3179 VDD.n1871 VDD.n1870 4.5005
R3180 VDD.n1803 VDD.n359 4.5005
R3181 VDD.n1685 VDD.n1684 4.5005
R3182 VDD.n1683 VDD.n1682 4.5005
R3183 VDD.n1620 VDD.n456 4.5005
R3184 VDD.n1526 VDD.n1525 4.5005
R3185 VDD.n1524 VDD.n1523 4.5005
R3186 VDD.n2301 VDD.n215 4.5005
R3187 VDD.n680 VDD.n679 4.5005
R3188 VDD.n2332 VDD.n2331 4.5005
R3189 VDD.n2219 VDD.n216 4.5005
R3190 VDD.n2152 VDD.n2151 4.5005
R3191 VDD.n2150 VDD.n2149 4.5005
R3192 VDD.n2058 VDD.n240 4.5005
R3193 VDD.n2002 VDD.n2001 4.5005
R3194 VDD.n2000 VDD.n1999 4.5005
R3195 VDD.n1896 VDD.n308 4.5005
R3196 VDD.n1838 VDD.n1837 4.5005
R3197 VDD.n1836 VDD.n1835 4.5005
R3198 VDD.n1710 VDD.n379 4.5005
R3199 VDD.n1644 VDD.n1643 4.5005
R3200 VDD.n1642 VDD.n1641 4.5005
R3201 VDD.n1551 VDD.n480 4.5005
R3202 VDD.n1483 VDD.n1482 4.5005
R3203 VDD.n2255 VDD.n2254 4.5005
R3204 VDD.n2253 VDD.n2252 4.5005
R3205 VDD.n772 VDD.n221 4.5005
R3206 VDD.n2083 VDD.n2082 4.5005
R3207 VDD.n2081 VDD.n2080 4.5005
R3208 VDD.n946 VDD.n252 4.5005
R3209 VDD.n1922 VDD.n1921 4.5005
R3210 VDD.n1920 VDD.n1919 4.5005
R3211 VDD.n1126 VDD.n319 4.5005
R3212 VDD.n1743 VDD.n1742 4.5005
R3213 VDD.n1741 VDD.n1740 4.5005
R3214 VDD.n1302 VDD.n406 4.5005
R3215 VDD.n1577 VDD.n1576 4.5005
R3216 VDD.n1575 VDD.n1574 4.5005
R3217 VDD.n1452 VDD.n499 4.5005
R3218 VDD.n145 VDD.n0 4.5005
R3219 VDD.n147 VDD.n146 4.5005
R3220 VDD.n148 VDD.n141 4.5005
R3221 VDD.n150 VDD.n149 4.5005
R3222 VDD.n151 VDD.n140 4.5005
R3223 VDD.n153 VDD.n152 4.5005
R3224 VDD.n155 VDD.n154 4.5005
R3225 VDD.n156 VDD.n138 4.5005
R3226 VDD.n158 VDD.n157 4.5005
R3227 VDD.n159 VDD.n137 4.5005
R3228 VDD.n161 VDD.n160 4.5005
R3229 VDD.n162 VDD.n136 4.5005
R3230 VDD.n164 VDD.n163 4.5005
R3231 VDD.n166 VDD.n165 4.5005
R3232 VDD.n167 VDD.n131 4.5005
R3233 VDD.n169 VDD.n168 4.5005
R3234 VDD.n170 VDD.n130 4.5005
R3235 VDD.n172 VDD.n171 4.5005
R3236 VDD.n173 VDD.n129 4.5005
R3237 VDD.n175 VDD.n174 4.5005
R3238 VDD.n100 VDD.n99 4.5005
R3239 VDD.n101 VDD.n14 4.5005
R3240 VDD.n103 VDD.n102 4.5005
R3241 VDD.n104 VDD.n13 4.5005
R3242 VDD.n106 VDD.n105 4.5005
R3243 VDD.n107 VDD.n1 4.5005
R3244 VDD.n1438 VDD.t14 4.46351
R3245 VDD.n1441 VDD.t694 4.46351
R3246 VDD.n1570 VDD.t3052 4.46351
R3247 VDD.n1569 VDD.t795 4.46351
R3248 VDD.n1553 VDD.t616 4.46351
R3249 VDD.n1550 VDD.t3221 4.46351
R3250 VDD.n1309 VDD.t3231 4.46351
R3251 VDD.n1307 VDD.t3472 4.46351
R3252 VDD.n1296 VDD.t806 4.46351
R3253 VDD.n1294 VDD.t2820 4.46351
R3254 VDD.n1299 VDD.t3609 4.46351
R3255 VDD.n1300 VDD.t785 4.46351
R3256 VDD.n1301 VDD.t3480 4.46351
R3257 VDD.n1303 VDD.t1809 4.46351
R3258 VDD.n1750 VDD.t3095 4.46351
R3259 VDD.n1752 VDD.t1037 4.46351
R3260 VDD.n1116 VDD.t4116 4.46351
R3261 VDD.n1114 VDD.t3756 4.46351
R3262 VDD.n1843 VDD.t3097 4.46351
R3263 VDD.n1911 VDD.t4110 4.46351
R3264 VDD.n1910 VDD.t1772 4.46351
R3265 VDD.n1909 VDD.t1067 4.46351
R3266 VDD.n1908 VDD.t3859 4.46351
R3267 VDD.n1885 VDD.t2425 4.46351
R3268 VDD.n1930 VDD.t10 4.46351
R3269 VDD.n1931 VDD.t896 4.46351
R3270 VDD.n2143 VDD.t16 4.46351
R3271 VDD.n2141 VDD.t3599 4.46351
R3272 VDD.n2133 VDD.t4108 4.46351
R3273 VDD.n2131 VDD.t2239 4.46351
R3274 VDD.n2166 VDD.t4058 4.46351
R3275 VDD.n2167 VDD.t635 4.46351
R3276 VDD.n2169 VDD.t4113 4.46351
R3277 VDD.n2170 VDD.t2545 4.46351
R3278 VDD.n650 VDD.t3808 4.39052
R3279 VDD.n621 VDD.t58 4.38377
R3280 VDD.n1497 VDD.t1701 4.36426
R3281 VDD.n1739 VDD.t2994 4.36426
R3282 VDD.n1737 VDD.t2327 4.36426
R3283 VDD.n1709 VDD.t4027 4.36426
R3284 VDD.n1726 VDD.t3699 4.36426
R3285 VDD.n1847 VDD.t1083 4.36426
R3286 VDD.n1858 VDD.t4275 4.36426
R3287 VDD.n1104 VDD.t849 4.36426
R3288 VDD.n1991 VDD.t789 4.36426
R3289 VDD.n307 VDD.t1835 4.36426
R3290 VDD.n2118 VDD.t2417 4.36426
R3291 VDD.n2165 VDD.t2465 4.36426
R3292 VDD.n2172 VDD.t3717 4.36426
R3293 VDD.n231 VDD.t2234 4.36426
R3294 VDD.n623 VDD.t1825 4.36035
R3295 VDD.n634 VDD.t2582 4.36035
R3296 VDD.n1385 VDD.t2230 4.36035
R3297 VDD.n1385 VDD.t2024 4.36035
R3298 VDD.n1377 VDD.t2664 4.36035
R3299 VDD.n1373 VDD.t3771 4.36035
R3300 VDD.n1414 VDD.t3197 4.36035
R3301 VDD.n1409 VDD.t3298 4.36035
R3302 VDD.n1411 VDD.t2961 4.36035
R3303 VDD.n1376 VDD.t3545 4.36035
R3304 VDD.n1378 VDD.t2957 4.36035
R3305 VDD.n1379 VDD.t913 4.36035
R3306 VDD.n1381 VDD.t2171 4.36035
R3307 VDD.n1382 VDD.t2443 4.36035
R3308 VDD.n1384 VDD.t3401 4.36035
R3309 VDD.n1339 VDD.t2658 4.36035
R3310 VDD.n1339 VDD.t4162 4.36035
R3311 VDD.n1338 VDD.t1503 4.36035
R3312 VDD.n1338 VDD.t2325 4.36035
R3313 VDD.n1337 VDD.t2441 4.36035
R3314 VDD.n1337 VDD.t4263 4.36035
R3315 VDD.n1336 VDD.t1488 4.36035
R3316 VDD.n1336 VDD.t1159 4.36035
R3317 VDD.n1335 VDD.t2195 4.36035
R3318 VDD.n1335 VDD.t2365 4.36035
R3319 VDD.n1334 VDD.t3038 4.36035
R3320 VDD.n1334 VDD.t3656 4.36035
R3321 VDD.n1333 VDD.t2549 4.36035
R3322 VDD.n1333 VDD.t3533 4.36035
R3323 VDD.n1368 VDD.t3069 4.36035
R3324 VDD.n1368 VDD.t3268 4.36035
R3325 VDD.n1364 VDD.t3294 4.36035
R3326 VDD.n1359 VDD.t4136 4.36035
R3327 VDD.n1365 VDD.t3912 4.36035
R3328 VDD.n1367 VDD.t3296 4.36035
R3329 VDD.n1370 VDD.t1805 4.36035
R3330 VDD.n1260 VDD.t2760 4.36035
R3331 VDD.n1258 VDD.t3579 4.36035
R3332 VDD.n1256 VDD.t2781 4.36035
R3333 VDD.n1254 VDD.t983 4.36035
R3334 VDD.n1252 VDD.t1215 4.36035
R3335 VDD.n1250 VDD.t2026 4.36035
R3336 VDD.n1248 VDD.t4289 4.36035
R3337 VDD.n1327 VDD.t2818 4.36035
R3338 VDD.n1325 VDD.t2570 4.36035
R3339 VDD.n1323 VDD.t2783 4.36035
R3340 VDD.n1321 VDD.t2482 4.36035
R3341 VDD.n1319 VDD.t2680 4.36035
R3342 VDD.n1317 VDD.t1436 4.36035
R3343 VDD.n1315 VDD.t3304 4.36035
R3344 VDD.n1313 VDD.t1021 4.36035
R3345 VDD.n1311 VDD.t2756 4.36035
R3346 VDD.n1306 VDD.t1161 4.36035
R3347 VDD.n1308 VDD.t2947 4.36035
R3348 VDD.n1310 VDD.t3317 4.36035
R3349 VDD.n1314 VDD.t942 4.36035
R3350 VDD.n1316 VDD.t3086 4.36035
R3351 VDD.n1318 VDD.t2891 4.36035
R3352 VDD.n1320 VDD.t3514 4.36035
R3353 VDD.n1322 VDD.t1888 4.36035
R3354 VDD.n1324 VDD.t2150 4.36035
R3355 VDD.n1326 VDD.t3334 4.36035
R3356 VDD.n1328 VDD.t3321 4.36035
R3357 VDD.n1330 VDD.t2308 4.36035
R3358 VDD.n1249 VDD.t2682 4.36035
R3359 VDD.n1251 VDD.t1581 4.36035
R3360 VDD.n1253 VDD.t3465 4.36035
R3361 VDD.n1255 VDD.t3837 4.36035
R3362 VDD.n1257 VDD.t3046 4.36035
R3363 VDD.n1259 VDD.t3207 4.36035
R3364 VDD.n1261 VDD.t4295 4.36035
R3365 VDD.n1219 VDD.t2152 4.36035
R3366 VDD.n1217 VDD.t3748 4.36035
R3367 VDD.n1215 VDD.t2130 4.36035
R3368 VDD.n1213 VDD.t2364 4.36035
R3369 VDD.n1211 VDD.t3822 4.36035
R3370 VDD.n1209 VDD.t3916 4.36035
R3371 VDD.n1207 VDD.t3847 4.36035
R3372 VDD.n1243 VDD.t3532 4.36035
R3373 VDD.n1241 VDD.t3418 4.36035
R3374 VDD.n1239 VDD.t3874 4.36035
R3375 VDD.n1237 VDD.t3914 4.36035
R3376 VDD.n1235 VDD.t2674 4.36035
R3377 VDD.n1233 VDD.t2072 4.36035
R3378 VDD.n1231 VDD.t1538 4.36035
R3379 VDD.n1229 VDD.t1117 4.36035
R3380 VDD.n1227 VDD.t3615 4.36035
R3381 VDD.n1225 VDD.t3530 4.36035
R3382 VDD.n1225 VDD.t1456 4.36035
R3383 VDD.n1224 VDD.t1924 4.36035
R3384 VDD.n1224 VDD.t1547 4.36035
R3385 VDD.n1223 VDD.t2229 4.36035
R3386 VDD.n1223 VDD.t3208 4.36035
R3387 VDD.n1222 VDD.t2795 4.36035
R3388 VDD.n1222 VDD.t2802 4.36035
R3389 VDD.n407 VDD.t4034 4.36035
R3390 VDD.n1221 VDD.t3611 4.36035
R3391 VDD.n1228 VDD.t2559 4.36035
R3392 VDD.n1230 VDD.t2935 4.36035
R3393 VDD.n1232 VDD.t1432 4.36035
R3394 VDD.n1234 VDD.t2540 4.36035
R3395 VDD.n1236 VDD.t3794 4.36035
R3396 VDD.n1238 VDD.t2710 4.36035
R3397 VDD.n1240 VDD.t958 4.36035
R3398 VDD.n1242 VDD.t1501 4.36035
R3399 VDD.n1245 VDD.t894 4.36035
R3400 VDD.n1208 VDD.t3203 4.36035
R3401 VDD.n1210 VDD.t1987 4.36035
R3402 VDD.n1212 VDD.t2889 4.36035
R3403 VDD.n1214 VDD.t2135 4.36035
R3404 VDD.n1216 VDD.t2392 4.36035
R3405 VDD.n1218 VDD.t2183 4.36035
R3406 VDD.n1220 VDD.t2250 4.36035
R3407 VDD.n1173 VDD.t3790 4.36035
R3408 VDD.n1171 VDD.t4212 4.36035
R3409 VDD.n1169 VDD.t1474 4.36035
R3410 VDD.n1167 VDD.t4267 4.36035
R3411 VDD.n1165 VDD.t1208 4.36035
R3412 VDD.n1163 VDD.t3251 4.36035
R3413 VDD.n1161 VDD.t3133 4.36035
R3414 VDD.n1201 VDD.t3970 4.36035
R3415 VDD.n1199 VDD.t3557 4.36035
R3416 VDD.n1197 VDD.t3550 4.36035
R3417 VDD.n1195 VDD.t1631 4.36035
R3418 VDD.n1193 VDD.t2124 4.36035
R3419 VDD.n1191 VDD.t2702 4.36035
R3420 VDD.n1189 VDD.t991 4.36035
R3421 VDD.n1187 VDD.t3765 4.36035
R3422 VDD.n1185 VDD.t970 4.36035
R3423 VDD.n1183 VDD.t3946 4.36035
R3424 VDD.n1744 VDD.t1452 4.36035
R3425 VDD.n1746 VDD.t2574 4.36035
R3426 VDD.n1181 VDD.t2648 4.36035
R3427 VDD.n1182 VDD.t2179 4.36035
R3428 VDD.n1184 VDD.t3010 4.36035
R3429 VDD.n1188 VDD.t2107 4.36035
R3430 VDD.n1190 VDD.t2553 4.36035
R3431 VDD.n1192 VDD.t1300 4.36035
R3432 VDD.n1194 VDD.t2419 4.36035
R3433 VDD.n1196 VDD.t3135 4.36035
R3434 VDD.n1198 VDD.t2447 4.36035
R3435 VDD.n1200 VDD.t3884 4.36035
R3436 VDD.n1202 VDD.t3099 4.36035
R3437 VDD.n1204 VDD.t3002 4.36035
R3438 VDD.n1162 VDD.t2396 4.36035
R3439 VDD.n1164 VDD.t2484 4.36035
R3440 VDD.n1166 VDD.t2014 4.36035
R3441 VDD.n1168 VDD.t1355 4.36035
R3442 VDD.n1170 VDD.t3247 4.36035
R3443 VDD.n1172 VDD.t3174 4.36035
R3444 VDD.n1174 VDD.t4291 4.36035
R3445 VDD.n1087 VDD.t1627 4.36035
R3446 VDD.n1085 VDD.t2913 4.36035
R3447 VDD.n1083 VDD.t2032 4.36035
R3448 VDD.n1081 VDD.t1913 4.36035
R3449 VDD.n1079 VDD.t1923 4.36035
R3450 VDD.n1077 VDD.t3940 4.36035
R3451 VDD.n1075 VDD.t1723 4.36035
R3452 VDD.n1156 VDD.t2899 4.36035
R3453 VDD.n1154 VDD.t4021 4.36035
R3454 VDD.n1152 VDD.t1993 4.36035
R3455 VDD.n1150 VDD.t1340 4.36035
R3456 VDD.n1148 VDD.t2322 4.36035
R3457 VDD.n1146 VDD.t2943 4.36035
R3458 VDD.n1144 VDD.t3399 4.36035
R3459 VDD.n1142 VDD.t3071 4.36035
R3460 VDD.n1140 VDD.t4182 4.36035
R3461 VDD.n1138 VDD.t2678 4.36035
R3462 VDD.n1136 VDD.t3525 4.36035
R3463 VDD.n1134 VDD.t3968 4.36035
R3464 VDD.n1132 VDD.t3130 4.36035
R3465 VDD.n1130 VDD.t2445 4.36035
R3466 VDD.n1128 VDD.t1524 4.36035
R3467 VDD.n1125 VDD.t3407 4.36035
R3468 VDD.n1123 VDD.t2113 4.36035
R3469 VDD.n1119 VDD.t2394 4.36035
R3470 VDD.n1120 VDD.t1244 4.36035
R3471 VDD.n1122 VDD.t4067 4.36035
R3472 VDD.n1124 VDD.t1236 4.36035
R3473 VDD.n1127 VDD.t2270 4.36035
R3474 VDD.n1129 VDD.t1359 4.36035
R3475 VDD.n1131 VDD.t4073 4.36035
R3476 VDD.n1133 VDD.t2875 4.36035
R3477 VDD.n1135 VDD.t2791 4.36035
R3478 VDD.n1137 VDD.t2666 4.36035
R3479 VDD.n1141 VDD.t3812 4.36035
R3480 VDD.n1143 VDD.t1841 4.36035
R3481 VDD.n1145 VDD.t4054 4.36035
R3482 VDD.n1147 VDD.t4106 4.36035
R3483 VDD.n1149 VDD.t4184 4.36035
R3484 VDD.n1151 VDD.t2037 4.36035
R3485 VDD.n1153 VDD.t1858 4.36035
R3486 VDD.n1155 VDD.t1444 4.36035
R3487 VDD.n1158 VDD.t968 4.36035
R3488 VDD.n1076 VDD.t1412 4.36035
R3489 VDD.n1078 VDD.t3454 4.36035
R3490 VDD.n1080 VDD.t3118 4.36035
R3491 VDD.n1082 VDD.t3342 4.36035
R3492 VDD.n1084 VDD.t2381 4.36035
R3493 VDD.n1086 VDD.t2292 4.36035
R3494 VDD.n1088 VDD.t2523 4.36035
R3495 VDD.n1040 VDD.t3804 4.36035
R3496 VDD.n1038 VDD.t2120 4.36035
R3497 VDD.n1036 VDD.t2028 4.36035
R3498 VDD.n1034 VDD.t3249 4.36035
R3499 VDD.n1032 VDD.t2869 4.36035
R3500 VDD.n1030 VDD.t1292 4.36035
R3501 VDD.n1028 VDD.t3577 4.36035
R3502 VDD.n1070 VDD.t2331 4.36035
R3503 VDD.n1068 VDD.t3008 4.36035
R3504 VDD.n1066 VDD.t3683 4.36035
R3505 VDD.n1064 VDD.t3109 4.36035
R3506 VDD.n1062 VDD.t976 4.36035
R3507 VDD.n1060 VDD.t2360 4.36035
R3508 VDD.n1058 VDD.t3143 4.36035
R3509 VDD.n1056 VDD.t4069 4.36035
R3510 VDD.n1054 VDD.t1131 4.36035
R3511 VDD.n1051 VDD.t3523 4.36035
R3512 VDD.n1049 VDD.t2300 4.36035
R3513 VDD.n1047 VDD.t3854 4.36035
R3514 VDD.n1045 VDD.t1416 4.36035
R3515 VDD.n1043 VDD.t1911 4.36035
R3516 VDD.n320 VDD.t1234 4.36035
R3517 VDD.n1917 VDD.t2591 4.36035
R3518 VDD.n1915 VDD.t3312 4.36035
R3519 VDD.n1912 VDD.t2754 4.36035
R3520 VDD.n1914 VDD.t2371 4.36035
R3521 VDD.n1916 VDD.t2810 4.36035
R3522 VDD.n1918 VDD.t3385 4.36035
R3523 VDD.n1042 VDD.t4198 4.36035
R3524 VDD.n1044 VDD.t3886 4.36035
R3525 VDD.n1046 VDD.t3263 4.36035
R3526 VDD.n1048 VDD.t3635 4.36035
R3527 VDD.n1050 VDD.t2547 4.36035
R3528 VDD.n1052 VDD.t2128 4.36035
R3529 VDD.n1055 VDD.t3752 4.36035
R3530 VDD.n1057 VDD.t2660 4.36035
R3531 VDD.n1059 VDD.t1410 4.36035
R3532 VDD.n1061 VDD.t3354 4.36035
R3533 VDD.n1063 VDD.t3516 4.36035
R3534 VDD.n1065 VDD.t3155 4.36035
R3535 VDD.n1067 VDD.t2676 4.36035
R3536 VDD.n1069 VDD.t1866 4.36035
R3537 VDD.n1072 VDD.t2584 4.36035
R3538 VDD.n1029 VDD.t4041 4.36035
R3539 VDD.n1031 VDD.t3568 4.36035
R3540 VDD.n1033 VDD.t999 4.36035
R3541 VDD.n1035 VDD.t4277 4.36035
R3542 VDD.n1037 VDD.t1915 4.36035
R3543 VDD.n1039 VDD.t3800 4.36035
R3544 VDD.n1041 VDD.t4283 4.36035
R3545 VDD.n993 VDD.t3746 4.36035
R3546 VDD.n991 VDD.t2963 4.36035
R3547 VDD.n989 VDD.t2871 4.36035
R3548 VDD.n987 VDD.t1511 4.36035
R3549 VDD.n985 VDD.t2039 4.36035
R3550 VDD.n983 VDD.t3894 4.36035
R3551 VDD.n981 VDD.t1629 4.36035
R3552 VDD.n1023 VDD.t4039 4.36035
R3553 VDD.n1021 VDD.t2369 4.36035
R3554 VDD.n1019 VDD.t2252 4.36035
R3555 VDD.n1017 VDD.t2254 4.36035
R3556 VDD.n1015 VDD.t1683 4.36035
R3557 VDD.n1013 VDD.t2861 4.36035
R3558 VDD.n1011 VDD.t1232 4.36035
R3559 VDD.n1009 VDD.t3280 4.36035
R3560 VDD.n1007 VDD.t1440 4.36035
R3561 VDD.n1004 VDD.t1801 4.36035
R3562 VDD.n1002 VDD.t3575 4.36035
R3563 VDD.n1000 VDD.t1813 4.36035
R3564 VDD.n998 VDD.t2102 4.36035
R3565 VDD.n996 VDD.t3088 4.36035
R3566 VDD.n318 VDD.t3987 4.36035
R3567 VDD.n1924 VDD.t2808 4.36035
R3568 VDD.n1926 VDD.t1811 4.36035
R3569 VDD.n1984 VDD.t2143 4.36035
R3570 VDD.n1929 VDD.t1133 4.36035
R3571 VDD.n1927 VDD.t3205 4.36035
R3572 VDD.n1925 VDD.t3587 4.36035
R3573 VDD.n1923 VDD.t1719 4.36035
R3574 VDD.n995 VDD.t2451 4.36035
R3575 VDD.n997 VDD.t2278 4.36035
R3576 VDD.n999 VDD.t4200 4.36035
R3577 VDD.n1001 VDD.t3573 4.36035
R3578 VDD.n1003 VDD.t2758 4.36035
R3579 VDD.n1005 VDD.t2494 4.36035
R3580 VDD.n1008 VDD.t3687 4.36035
R3581 VDD.n1010 VDD.t2490 4.36035
R3582 VDD.n1012 VDD.t4097 4.36035
R3583 VDD.n1014 VDD.t4043 4.36035
R3584 VDD.n1016 VDD.t3950 4.36035
R3585 VDD.n1018 VDD.t2670 4.36035
R3586 VDD.n1020 VDD.t2362 4.36035
R3587 VDD.n1022 VDD.t3199 4.36035
R3588 VDD.n1025 VDD.t2775 4.36035
R3589 VDD.n982 VDD.t978 4.36035
R3590 VDD.n984 VDD.t2668 4.36035
R3591 VDD.n986 VDD.t2215 4.36035
R3592 VDD.n988 VDD.t2897 4.36035
R3593 VDD.n990 VDD.t2730 4.36035
R3594 VDD.n992 VDD.t1790 4.36035
R3595 VDD.n994 VDD.t2799 4.36035
R3596 VDD.n913 VDD.t3592 4.36035
R3597 VDD.n911 VDD.t1135 4.36035
R3598 VDD.n909 VDD.t3075 4.36035
R3599 VDD.n907 VDD.t1583 4.36035
R3600 VDD.n905 VDD.t1139 4.36035
R3601 VDD.n903 VDD.t2726 4.36035
R3602 VDD.n901 VDD.t3082 4.36035
R3603 VDD.n976 VDD.t3942 4.36035
R3604 VDD.n974 VDD.t3319 4.36035
R3605 VDD.n972 VDD.t2844 4.36035
R3606 VDD.n970 VDD.t1213 4.36035
R3607 VDD.n968 VDD.t3989 4.36035
R3608 VDD.n966 VDD.t1708 4.36035
R3609 VDD.n964 VDD.t3839 4.36035
R3610 VDD.n962 VDD.t3239 4.36035
R3611 VDD.n960 VDD.t3044 4.36035
R3612 VDD.n958 VDD.t2708 4.36035
R3613 VDD.n956 VDD.t4239 4.36035
R3614 VDD.n954 VDD.t2824 4.36035
R3615 VDD.n952 VDD.t2302 4.36035
R3616 VDD.n950 VDD.t3188 4.36035
R3617 VDD.n948 VDD.t3291 4.36035
R3618 VDD.n945 VDD.t1731 4.36035
R3619 VDD.n943 VDD.t2836 4.36035
R3620 VDD.n939 VDD.t2030 4.36035
R3621 VDD.n937 VDD.t3370 4.36035
R3622 VDD.n935 VDD.t1985 4.36035
R3623 VDD.n933 VDD.t2555 4.36035
R3624 VDD.n2004 VDD.t4301 4.36035
R3625 VDD.n930 VDD.t2433 4.36035
R3626 VDD.n931 VDD.t2296 4.36035
R3627 VDD.n932 VDD.t3016 4.36035
R3628 VDD.n934 VDD.t1480 4.36035
R3629 VDD.n936 VDD.t1778 4.36035
R3630 VDD.n938 VDD.t2062 4.36035
R3631 VDD.n940 VDD.t3458 4.36035
R3632 VDD.n942 VDD.t3685 4.36035
R3633 VDD.n944 VDD.t985 4.36035
R3634 VDD.n947 VDD.t4233 4.36035
R3635 VDD.n949 VDD.t2085 4.36035
R3636 VDD.n951 VDD.t3422 4.36035
R3637 VDD.n953 VDD.t1890 4.36035
R3638 VDD.n955 VDD.t3833 4.36035
R3639 VDD.n957 VDD.t2202 4.36035
R3640 VDD.n961 VDD.t2093 4.36035
R3641 VDD.n963 VDD.t3163 4.36035
R3642 VDD.n965 VDD.t1938 4.36035
R3643 VDD.n967 VDD.t1536 4.36035
R3644 VDD.n969 VDD.t1424 4.36035
R3645 VDD.n971 VDD.t2421 4.36035
R3646 VDD.n973 VDD.t3948 4.36035
R3647 VDD.n975 VDD.t1621 4.36035
R3648 VDD.n978 VDD.t2941 4.36035
R3649 VDD.n902 VDD.t4214 4.36035
R3650 VDD.n904 VDD.t899 4.36035
R3651 VDD.n906 VDD.t4202 4.36035
R3652 VDD.n908 VDD.t2801 4.36035
R3653 VDD.n910 VDD.t1482 4.36035
R3654 VDD.n912 VDD.t4208 4.36035
R3655 VDD.n914 VDD.t3420 4.36035
R3656 VDD.n866 VDD.t1740 4.36035
R3657 VDD.n864 VDD.t3641 4.36035
R3658 VDD.n862 VDD.t3924 4.36035
R3659 VDD.n860 VDD.t1260 4.36035
R3660 VDD.n858 VDD.t2561 4.36035
R3661 VDD.n856 VDD.t3666 4.36035
R3662 VDD.n854 VDD.t4228 4.36035
R3663 VDD.n896 VDD.t2126 4.36035
R3664 VDD.n894 VDD.t3382 4.36035
R3665 VDD.n892 VDD.t3689 4.36035
R3666 VDD.n890 VDD.t3537 4.36035
R3667 VDD.n888 VDD.t2722 4.36035
R3668 VDD.n886 VDD.t3452 4.36035
R3669 VDD.n884 VDD.t3346 4.36035
R3670 VDD.n882 VDD.t3092 4.36035
R3671 VDD.n880 VDD.t2527 4.36035
R3672 VDD.n877 VDD.t1680 4.36035
R3673 VDD.n875 VDD.t3977 4.36035
R3674 VDD.n873 VDD.t966 4.36035
R3675 VDD.n871 VDD.t3930 4.36035
R3676 VDD.n869 VDD.t4000 4.36035
R3677 VDD.n253 VDD.t1733 4.36035
R3678 VDD.n2078 VDD.t1738 4.36035
R3679 VDD.n2076 VDD.t3137 4.36035
R3680 VDD.n2073 VDD.t4137 4.36035
R3681 VDD.n2073 VDD.t2324 4.36035
R3682 VDD.n2072 VDD.t2876 4.36035
R3683 VDD.n2072 VDD.t2267 4.36035
R3684 VDD.n2071 VDD.t3408 4.36035
R3685 VDD.n2071 VDD.t2148 4.36035
R3686 VDD.n2070 VDD.t1369 4.36035
R3687 VDD.n2070 VDD.t3258 4.36035
R3688 VDD.n2069 VDD.t1420 4.36035
R3689 VDD.n2069 VDD.t2646 4.36035
R3690 VDD.n2065 VDD.t2728 4.36035
R3691 VDD.n2067 VDD.t4079 4.36035
R3692 VDD.n2068 VDD.t4140 4.36035
R3693 VDD.n2075 VDD.t3627 4.36035
R3694 VDD.n2077 VDD.t2521 4.36035
R3695 VDD.n2079 VDD.t2641 4.36035
R3696 VDD.n868 VDD.t3253 4.36035
R3697 VDD.n870 VDD.t3378 4.36035
R3698 VDD.n872 VDD.t3529 4.36035
R3699 VDD.n874 VDD.t940 4.36035
R3700 VDD.n876 VDD.t1196 4.36035
R3701 VDD.n878 VDD.t1371 4.36035
R3702 VDD.n881 VDD.t2173 4.36035
R3703 VDD.n883 VDD.t1252 4.36035
R3704 VDD.n885 VDD.t1298 4.36035
R3705 VDD.n887 VDD.t2643 4.36035
R3706 VDD.n889 VDD.t4012 4.36035
R3707 VDD.n891 VDD.t1229 4.36035
R3708 VDD.n893 VDD.t1246 4.36035
R3709 VDD.n895 VDD.t4168 4.36035
R3710 VDD.n898 VDD.t2316 4.36035
R3711 VDD.n855 VDD.t3113 4.36035
R3712 VDD.n857 VDD.t1227 4.36035
R3713 VDD.n859 VDD.t4172 4.36035
R3714 VDD.n861 VDD.t4178 4.36035
R3715 VDD.n863 VDD.t2158 4.36035
R3716 VDD.n865 VDD.t3470 4.36035
R3717 VDD.n867 VDD.t3050 4.36035
R3718 VDD.n819 VDD.t2830 4.36035
R3719 VDD.n817 VDD.t2662 4.36035
R3720 VDD.n815 VDD.t4287 4.36035
R3721 VDD.n813 VDD.t2903 4.36035
R3722 VDD.n811 VDD.t3103 4.36035
R3723 VDD.n809 VDD.t2399 4.36035
R3724 VDD.n807 VDD.t2304 4.36035
R3725 VDD.n849 VDD.t3237 4.36035
R3726 VDD.n847 VDD.t1633 4.36035
R3727 VDD.n845 VDD.t1685 4.36035
R3728 VDD.n843 VDD.t3843 4.36035
R3729 VDD.n841 VDD.t3004 4.36035
R3730 VDD.n839 VDD.t3278 4.36035
R3731 VDD.n837 VDD.t1803 4.36035
R3732 VDD.n835 VDD.t2901 4.36035
R3733 VDD.n833 VDD.t3784 4.36035
R3734 VDD.n830 VDD.t2477 4.36035
R3735 VDD.n828 VDD.t4219 4.36035
R3736 VDD.n826 VDD.t3655 4.36035
R3737 VDD.n824 VDD.t3719 4.36035
R3738 VDD.n822 VDD.t2403 4.36035
R3739 VDD.n251 VDD.t2463 4.36035
R3740 VDD.n2085 VDD.t3014 4.36035
R3741 VDD.n2087 VDD.t1191 4.36035
R3742 VDD.n2090 VDD.t989 4.36035
R3743 VDD.n2090 VDD.t1394 4.36035
R3744 VDD.n2091 VDD.t4050 4.36035
R3745 VDD.n2091 VDD.t2777 4.36035
R3746 VDD.n2092 VDD.t2367 4.36035
R3747 VDD.n2092 VDD.t3763 4.36035
R3748 VDD.n2093 VDD.t954 4.36035
R3749 VDD.n2093 VDD.t1448 4.36035
R3750 VDD.n2094 VDD.t1839 4.36035
R3751 VDD.n2094 VDD.t1202 4.36035
R3752 VDD.n2095 VDD.t1681 4.36035
R3753 VDD.n2095 VDD.t1329 4.36035
R3754 VDD.n2096 VDD.t2386 4.36035
R3755 VDD.n2096 VDD.t3681 4.36035
R3756 VDD.n2097 VDD.t3992 4.36035
R3757 VDD.n2097 VDD.t3145 4.36035
R3758 VDD.n2098 VDD.t2720 4.36035
R3759 VDD.n2118 VDD.t2998 4.36035
R3760 VDD.n2117 VDD.t4138 4.36035
R3761 VDD.n2117 VDD.t1219 4.36035
R3762 VDD.n2116 VDD.t1788 4.36035
R3763 VDD.n2116 VDD.t4215 4.36035
R3764 VDD.n2120 VDD.t1792 4.36035
R3765 VDD.n2088 VDD.t3645 4.36035
R3766 VDD.n2086 VDD.t4159 4.36035
R3767 VDD.n2084 VDD.t4293 4.36035
R3768 VDD.n821 VDD.t3478 4.36035
R3769 VDD.n823 VDD.t972 4.36035
R3770 VDD.n825 VDD.t4170 4.36035
R3771 VDD.n827 VDD.t2043 4.36035
R3772 VDD.n829 VDD.t1991 4.36035
R3773 VDD.n831 VDD.t3153 4.36035
R3774 VDD.n834 VDD.t3426 4.36035
R3775 VDD.n836 VDD.t3006 4.36035
R3776 VDD.n838 VDD.t1351 4.36035
R3777 VDD.n840 VDD.t2955 4.36035
R3778 VDD.n842 VDD.t1983 4.36035
R3779 VDD.n844 VDD.t4102 4.36035
R3780 VDD.n846 VDD.t2840 4.36035
R3781 VDD.n848 VDD.t3882 4.36035
R3782 VDD.n851 VDD.t3157 4.36035
R3783 VDD.n808 VDD.t2449 4.36035
R3784 VDD.n810 VDD.t4077 4.36035
R3785 VDD.n812 VDD.t1100 4.36035
R3786 VDD.n814 VDD.t4281 4.36035
R3787 VDD.n816 VDD.t2160 4.36035
R3788 VDD.n818 VDD.t2210 4.36035
R3789 VDD.n820 VDD.t2008 4.36035
R3790 VDD.n740 VDD.t3424 4.36035
R3791 VDD.n738 VDD.t1333 4.36035
R3792 VDD.n736 VDD.t3964 4.36035
R3793 VDD.n734 VDD.t1617 4.36035
R3794 VDD.n732 VDD.t3996 4.36035
R3795 VDD.n730 VDD.t3042 4.36035
R3796 VDD.n728 VDD.t4226 4.36035
R3797 VDD.n802 VDD.t2276 4.36035
R3798 VDD.n800 VDD.t1762 4.36035
R3799 VDD.n798 VDD.t1290 4.36035
R3800 VDD.n796 VDD.t2945 4.36035
R3801 VDD.n794 VDD.t2298 4.36035
R3802 VDD.n792 VDD.t3179 4.36035
R3803 VDD.n790 VDD.t3637 4.36035
R3804 VDD.n788 VDD.t1180 4.36035
R3805 VDD.n786 VDD.t4273 4.36035
R3806 VDD.n783 VDD.t2653 4.36035
R3807 VDD.n781 VDD.t1422 4.36035
R3808 VDD.n779 VDD.t2486 4.36035
R3809 VDD.n777 VDD.t2992 4.36035
R3810 VDD.n775 VDD.t3972 4.36035
R3811 VDD.n773 VDD.t1725 4.36035
R3812 VDD.n770 VDD.t3428 4.36035
R3813 VDD.n768 VDD.t2873 4.36035
R3814 VDD.n765 VDD.t4104 4.36035
R3815 VDD.n763 VDD.t3159 4.36035
R3816 VDD.n761 VDD.t3672 4.36035
R3817 VDD.n759 VDD.t2576 4.36035
R3818 VDD.n757 VDD.t3436 4.36035
R3819 VDD.n755 VDD.t3267 4.36035
R3820 VDD.n753 VDD.t3585 4.36035
R3821 VDD.n751 VDD.t3035 4.36035
R3822 VDD.n749 VDD.t932 4.36035
R3823 VDD.n747 VDD.t915 4.36035
R3824 VDD.n745 VDD.t3241 4.36035
R3825 VDD.n743 VDD.t2816 4.36035
R3826 VDD.n239 VDD.t3101 4.36035
R3827 VDD.n2154 VDD.t4204 4.36035
R3828 VDD.n2156 VDD.t960 4.36035
R3829 VDD.n2162 VDD.t1770 4.36035
R3830 VDD.n231 VDD.t3559 4.36035
R3831 VDD.n2186 VDD.t2401 4.36035
R3832 VDD.n2184 VDD.t4269 4.36035
R3833 VDD.n2182 VDD.t1934 4.36035
R3834 VDD.n2180 VDD.t2885 4.36035
R3835 VDD.n2178 VDD.t4052 4.36035
R3836 VDD.n2176 VDD.t1663 4.36035
R3837 VDD.n2164 VDD.t3201 4.36035
R3838 VDD.n2163 VDD.t3270 4.36035
R3839 VDD.n2161 VDD.t1055 4.36035
R3840 VDD.n2159 VDD.t1338 4.36035
R3841 VDD.n2158 VDD.t3521 4.36035
R3842 VDD.n2157 VDD.t3680 4.36035
R3843 VDD.n2155 VDD.t3380 4.36035
R3844 VDD.n2153 VDD.t3938 4.36035
R3845 VDD.n742 VDD.t924 4.36035
R3846 VDD.n744 VDD.t3810 4.36035
R3847 VDD.n746 VDD.t1242 4.36035
R3848 VDD.n750 VDD.t3788 4.36035
R3849 VDD.n752 VDD.t3485 4.36035
R3850 VDD.n754 VDD.t2538 4.36035
R3851 VDD.n756 VDD.t3405 4.36035
R3852 VDD.n758 VDD.t1434 4.36035
R3853 VDD.n760 VDD.t3456 4.36035
R3854 VDD.n762 VDD.t1976 4.36035
R3855 VDD.n764 VDD.t2534 4.36035
R3856 VDD.n767 VDD.t1786 4.36035
R3857 VDD.n769 VDD.t2423 4.36035
R3858 VDD.n771 VDD.t2604 4.36035
R3859 VDD.n774 VDD.t2704 4.36035
R3860 VDD.n776 VDD.t3374 4.36035
R3861 VDD.n778 VDD.t1675 4.36035
R3862 VDD.n780 VDD.t1389 4.36035
R3863 VDD.n782 VDD.t2208 4.36035
R3864 VDD.n784 VDD.t1250 4.36035
R3865 VDD.n787 VDD.t2064 4.36035
R3866 VDD.n789 VDD.t1248 4.36035
R3867 VDD.n791 VDD.t934 4.36035
R3868 VDD.n793 VDD.t2373 4.36035
R3869 VDD.n795 VDD.t1833 4.36035
R3870 VDD.n797 VDD.t1418 4.36035
R3871 VDD.n799 VDD.t1098 4.36035
R3872 VDD.n801 VDD.t4151 4.36035
R3873 VDD.n804 VDD.t2256 4.36035
R3874 VDD.n729 VDD.t3111 4.36035
R3875 VDD.n731 VDD.t1225 4.36035
R3876 VDD.n733 VDD.t4157 4.36035
R3877 VDD.n735 VDD.t4164 4.36035
R3878 VDD.n737 VDD.t3643 4.36035
R3879 VDD.n739 VDD.t3806 4.36035
R3880 VDD.n741 VDD.t3450 4.36035
R3881 VDD.n693 VDD.t1472 4.36035
R3882 VDD.n691 VDD.t4271 4.36035
R3883 VDD.n689 VDD.t2832 4.36035
R3884 VDD.n687 VDD.t1558 4.36035
R3885 VDD.n685 VDD.t3120 4.36035
R3886 VDD.n683 VDD.t3372 4.36035
R3887 VDD.n681 VDD.t1187 4.36035
R3888 VDD.n723 VDD.t3868 4.36035
R3889 VDD.n721 VDD.t2959 4.36035
R3890 VDD.n719 VDD.t919 4.36035
R3891 VDD.n717 VDD.t928 4.36035
R3892 VDD.n715 VDD.t2980 4.36035
R3893 VDD.n713 VDD.t1344 4.36035
R3894 VDD.n711 VDD.t2580 4.36035
R3895 VDD.n709 VDD.t3918 4.36035
R3896 VDD.n707 VDD.t3440 4.36035
R3897 VDD.n704 VDD.t2405 4.36035
R3898 VDD.n702 VDD.t2834 4.36035
R3899 VDD.n700 VDD.t2967 4.36035
R3900 VDD.n698 VDD.t4144 4.36035
R3901 VDD.n696 VDD.t1150 4.36035
R3902 VDD.n222 VDD.t3368 4.36035
R3903 VDD.n2250 VDD.t2492 4.36035
R3904 VDD.n2248 VDD.t3936 4.36035
R3905 VDD.n2245 VDD.t2895 4.36035
R3906 VDD.n2243 VDD.t3828 4.36035
R3907 VDD.n2241 VDD.t1946 4.36035
R3908 VDD.n2239 VDD.t1635 4.36035
R3909 VDD.n2237 VDD.t3167 4.36035
R3910 VDD.n2235 VDD.t1899 4.36035
R3911 VDD.n2233 VDD.t1281 4.36035
R3912 VDD.n2231 VDD.t1104 4.36035
R3913 VDD.n2229 VDD.t3944 4.36035
R3914 VDD.n2226 VDD.t2272 4.36035
R3915 VDD.n2224 VDD.t2204 4.36035
R3916 VDD.n2222 VDD.t2154 4.36035
R3917 VDD.n2220 VDD.t2091 4.36035
R3918 VDD.n2217 VDD.t2221 4.36035
R3919 VDD.n2215 VDD.t2274 4.36035
R3920 VDD.n2213 VDD.t2265 4.36035
R3921 VDD.n2211 VDD.t2572 4.36035
R3922 VDD.n2207 VDD.t2797 4.36035
R3923 VDD.n2205 VDD.t2488 4.36035
R3924 VDD.n2203 VDD.t2116 4.36035
R3925 VDD.n2201 VDD.t3876 4.36035
R3926 VDD.n2198 VDD.t1143 4.36035
R3927 VDD.n2196 VDD.t2175 4.36035
R3928 VDD.n2194 VDD.t3539 4.36035
R3929 VDD.n2192 VDD.t3829 4.36035
R3930 VDD.n2192 VDD.t1585 4.36035
R3931 VDD.n229 VDD.t3209 4.36035
R3932 VDD.n229 VDD.t1608 4.36035
R3933 VDD.n228 VDD.t3555 4.36035
R3934 VDD.n228 VDD.t4032 4.36035
R3935 VDD.n227 VDD.t4229 4.36035
R3936 VDD.n227 VDD.t3336 4.36035
R3937 VDD.n226 VDD.t3344 4.36035
R3938 VDD.n226 VDD.t3562 4.36035
R3939 VDD.n225 VDD.t1240 4.36035
R3940 VDD.n225 VDD.t3852 4.36035
R3941 VDD.n224 VDD.t2114 4.36035
R3942 VDD.n224 VDD.t1610 4.36035
R3943 VDD.n223 VDD.t909 4.36035
R3944 VDD.n223 VDD.t3313 4.36035
R3945 VDD.n2195 VDD.t1970 4.36035
R3946 VDD.n2197 VDD.t1989 4.36035
R3947 VDD.n2199 VDD.t2458 4.36035
R3948 VDD.n2200 VDD.t1442 4.36035
R3949 VDD.n2202 VDD.t3302 4.36035
R3950 VDD.n2204 VDD.t4237 4.36035
R3951 VDD.n2206 VDD.t2838 4.36035
R3952 VDD.n2208 VDD.t2456 4.36035
R3953 VDD.n2210 VDD.t2511 4.36035
R3954 VDD.n2212 VDD.t3147 4.36035
R3955 VDD.n2214 VDD.t3170 4.36035
R3956 VDD.n2216 VDD.t2473 4.36035
R3957 VDD.n2218 VDD.t1576 4.36035
R3958 VDD.n2221 VDD.t3181 4.36035
R3959 VDD.n2223 VDD.t3315 4.36035
R3960 VDD.n2225 VDD.t1106 4.36035
R3961 VDD.n2227 VDD.t2469 4.36035
R3962 VDD.n2230 VDD.t2517 4.36035
R3963 VDD.n2232 VDD.t3172 4.36035
R3964 VDD.n2234 VDD.t875 4.36035
R3965 VDD.n2236 VDD.t3878 4.36035
R3966 VDD.n2238 VDD.t3779 4.36035
R3967 VDD.n2240 VDD.t905 4.36035
R3968 VDD.n2242 VDD.t3306 4.36035
R3969 VDD.n2244 VDD.t3831 4.36035
R3970 VDD.n2247 VDD.t2812 4.36035
R3971 VDD.n2249 VDD.t1794 4.36035
R3972 VDD.n2251 VDD.t1438 4.36035
R3973 VDD.n695 VDD.t3165 4.36035
R3974 VDD.n697 VDD.t2846 4.36035
R3975 VDD.n699 VDD.t3161 4.36035
R3976 VDD.n701 VDD.t2217 4.36035
R3977 VDD.n703 VDD.t1540 4.36035
R3978 VDD.n705 VDD.t1980 4.36035
R3979 VDD.n708 VDD.t1137 4.36035
R3980 VDD.n710 VDD.t3594 4.36035
R3981 VDD.n712 VDD.t3442 4.36035
R3982 VDD.n714 VDD.t1499 4.36035
R3983 VDD.n716 VDD.t936 4.36035
R3984 VDD.n718 VDD.t3713 4.36035
R3985 VDD.n720 VDD.t2415 4.36035
R3986 VDD.n722 VDD.t2850 4.36035
R3987 VDD.n725 VDD.t3709 4.36035
R3988 VDD.n682 VDD.t1322 4.36035
R3989 VDD.n684 VDD.t2822 4.36035
R3990 VDD.n686 VDD.t3674 4.36035
R3991 VDD.n688 VDD.t4006 4.36035
R3992 VDD.n690 VDD.t1901 4.36035
R3993 VDD.n692 VDD.t1346 4.36035
R3994 VDD.n694 VDD.t2865 4.36035
R3995 VDD.n648 VDD.t1560 4.36035
R3996 VDD.n646 VDD.t1516 4.36035
R3997 VDD.n644 VDD.t3397 4.36035
R3998 VDD.n642 VDD.t2598 4.36035
R3999 VDD.n640 VDD.t3890 4.36035
R4000 VDD.n638 VDD.t1148 4.36035
R4001 VDD.n677 VDD.t1294 4.36035
R4002 VDD.n677 VDD.t4296 4.36035
R4003 VDD.n676 VDD.t901 4.36035
R4004 VDD.n673 VDD.t1189 4.36035
R4005 VDD.n671 VDD.t3814 4.36035
R4006 VDD.n669 VDD.t2306 4.36035
R4007 VDD.n667 VDD.t3928 4.36035
R4008 VDD.n665 VDD.t4161 4.36035
R4009 VDD.n663 VDD.t950 4.36035
R4010 VDD.n661 VDD.t2156 4.36035
R4011 VDD.n659 VDD.t4016 4.36035
R4012 VDD.n657 VDD.t3564 4.36035
R4013 VDD.n657 VDD.t4017 4.36035
R4014 VDD.n656 VDD.t3168 4.36035
R4015 VDD.n656 VDD.t2045 4.36035
R4016 VDD.n655 VDD.t987 4.36035
R4017 VDD.n655 VDD.t3870 4.36035
R4018 VDD.n654 VDD.t4098 4.36035
R4019 VDD.n654 VDD.t2193 4.36035
R4020 VDD.n220 VDD.t3012 4.36035
R4021 VDD.n220 VDD.t3056 4.36035
R4022 VDD.n2256 VDD.t962 4.36035
R4023 VDD.n2256 VDD.t2243 4.36035
R4024 VDD.n2257 VDD.t3292 4.36035
R4025 VDD.n2257 VDD.t2779 4.36035
R4026 VDD.n2260 VDD.t2237 4.36035
R4027 VDD.n2262 VDD.t3036 4.36035
R4028 VDD.n2262 VDD.t2095 4.36035
R4029 VDD.n2263 VDD.t1003 4.36035
R4030 VDD.n2263 VDD.t3383 4.36035
R4031 VDD.n2264 VDD.t3468 4.36035
R4032 VDD.n2264 VDD.t1462 4.36035
R4033 VDD.n2265 VDD.t2087 4.36035
R4034 VDD.n2265 VDD.t3869 4.36035
R4035 VDD.n2266 VDD.t2248 4.36035
R4036 VDD.n2266 VDD.t2219 4.36035
R4037 VDD.n2267 VDD.t2856 4.36035
R4038 VDD.n2267 VDD.t2793 4.36035
R4039 VDD.n2268 VDD.t1163 4.36035
R4040 VDD.n2268 VDD.t2056 4.36035
R4041 VDD.n2269 VDD.t3724 4.36035
R4042 VDD.n2269 VDD.t2049 4.36035
R4043 VDD.n2270 VDD.t1402 4.36035
R4044 VDD.n2274 VDD.t3326 4.36035
R4045 VDD.n2272 VDD.t2167 4.36035
R4046 VDD.n217 VDD.t1864 4.36035
R4047 VDD.n2329 VDD.t2070 4.36035
R4048 VDD.n2327 VDD.t1406 4.36035
R4049 VDD.n2325 VDD.t4254 4.36035
R4050 VDD.n2323 VDD.t2996 4.36035
R4051 VDD.n2320 VDD.t4056 4.36035
R4052 VDD.n2318 VDD.t3352 4.36035
R4053 VDD.n2316 VDD.t1342 4.36035
R4054 VDD.n2314 VDD.t3387 4.36035
R4055 VDD.n2313 VDD.t3149 4.36035
R4056 VDD.n2311 VDD.t2771 4.36035
R4057 VDD.n2309 VDD.t2206 4.36035
R4058 VDD.n2307 VDD.t1217 4.36035
R4059 VDD.n2305 VDD.t2197 4.36035
R4060 VDD.n2303 VDD.t2586 4.36035
R4061 VDD.n2300 VDD.t4075 4.36035
R4062 VDD.n2298 VDD.t1206 4.36035
R4063 VDD.n2296 VDD.t3227 4.36035
R4064 VDD.n2294 VDD.t2939 4.36035
R4065 VDD.n2292 VDD.t1852 4.36035
R4066 VDD.n2290 VDD.t4100 4.36035
R4067 VDD.n2288 VDD.t3775 4.36035
R4068 VDD.n2302 VDD.t1764 4.36035
R4069 VDD.n2306 VDD.t4256 4.36035
R4070 VDD.n2308 VDD.t3998 4.36035
R4071 VDD.n2310 VDD.t4279 4.36035
R4072 VDD.n2312 VDD.t2018 4.36035
R4073 VDD.n2317 VDD.t4002 4.36035
R4074 VDD.n2322 VDD.t4004 4.36035
R4075 VDD.n2324 VDD.t2773 4.36035
R4076 VDD.n2326 VDD.t1170 4.36035
R4077 VDD.n2328 VDD.t1522 4.36035
R4078 VDD.n2330 VDD.t3272 4.36035
R4079 VDD.n2271 VDD.t4265 4.36035
R4080 VDD.n2273 VDD.t2379 4.36035
R4081 VDD.n2275 VDD.t2068 4.36035
R4082 VDD.n2258 VDD.t2047 4.36035
R4083 VDD.n660 VDD.t2645 4.36035
R4084 VDD.n662 VDD.t3566 4.36035
R4085 VDD.n664 VDD.t3726 4.36035
R4086 VDD.n666 VDD.t3979 4.36035
R4087 VDD.n668 VDD.t2318 4.36035
R4088 VDD.n670 VDD.t1619 4.36035
R4089 VDD.n672 VDD.t952 4.36035
R4090 VDD.n674 VDD.t3211 4.36035
R4091 VDD.n637 VDD.t4049 4.36035
R4092 VDD.n639 VDD.t3492 4.36035
R4093 VDD.n641 VDD.t2388 4.36035
R4094 VDD.n643 VDD.t3857 4.36035
R4095 VDD.n645 VDD.t1562 4.36035
R4096 VDD.n647 VDD.t1458 4.36035
R4097 VDD.n649 VDD.t3707 4.36035
R4098 VDD.n1439 VDD.n601 4.35924
R4099 VDD.n1406 VDD.n1393 4.35924
R4100 VDD.n1357 VDD.n1346 4.35924
R4101 VDD.n1312 VDD.n1262 4.35924
R4102 VDD.n1226 VDD.t3614 4.35924
R4103 VDD.n1186 VDD.n1175 4.35924
R4104 VDD.n1139 VDD.t4181 4.35924
R4105 VDD.n1053 VDD.t1130 4.35924
R4106 VDD.n1006 VDD.t1439 4.35924
R4107 VDD.n959 VDD.t3043 4.35924
R4108 VDD.n879 VDD.t2526 4.35924
R4109 VDD.n832 VDD.t3783 4.35924
R4110 VDD.n785 VDD.t4272 4.35924
R4111 VDD.n706 VDD.t3439 4.35924
R4112 VDD.n1508 VDD.n1507 4.35923
R4113 VDD.n1494 VDD.n566 4.35923
R4114 VDD.n1476 VDD.n576 4.35923
R4115 VDD.n1425 VDD.n610 4.35923
R4116 VDD.n1442 VDD.n600 4.35923
R4117 VDD.n1460 VDD.n586 4.35923
R4118 VDD.n1545 VDD.n517 4.35923
R4119 VDD.n1568 VDD.n502 4.35923
R4120 VDD.n1416 VDD.n1386 4.35923
R4121 VDD.n1633 VDD.n1598 4.35923
R4122 VDD.n1369 VDD.n1340 4.35923
R4123 VDD.n1580 VDD.n494 4.35923
R4124 VDD.n1654 VDD.n473 4.35923
R4125 VDD.n1329 VDD.t2307 4.35923
R4126 VDD.n1298 VDD.n1265 4.35923
R4127 VDD.n1699 VDD.n432 4.35923
R4128 VDD.n1244 VDD.t893 4.35923
R4129 VDD.n1735 VDD.n409 4.35923
R4130 VDD.n1824 VDD.n1776 4.35923
R4131 VDD.n1203 VDD.t3001 4.35923
R4132 VDD.n1748 VDD.n401 4.35923
R4133 VDD.n1845 VDD.n373 4.35923
R4134 VDD.n1157 VDD.t967 4.35923
R4135 VDD.n1121 VDD.n1089 4.35923
R4136 VDD.n1071 VDD.t2583 4.35923
R4137 VDD.n1913 VDD.t2370 4.35923
R4138 VDD.n1886 VDD.n334 4.35923
R4139 VDD.n1992 VDD.n1950 4.35923
R4140 VDD.n1024 VDD.t2774 4.35923
R4141 VDD.n1928 VDD.t3204 4.35923
R4142 VDD.n977 VDD.t2940 4.35923
R4143 VDD.n941 VDD.n915 4.35923
R4144 VDD.n2008 VDD.n303 4.35923
R4145 VDD.n2050 VDD.n262 4.35923
R4146 VDD.n897 VDD.t2315 4.35923
R4147 VDD.n2074 VDD.t3626 4.35923
R4148 VDD.n850 VDD.t3156 4.35923
R4149 VDD.n2089 VDD.t3644 4.35923
R4150 VDD.n2140 VDD.n2104 4.35923
R4151 VDD.n803 VDD.t2255 4.35923
R4152 VDD.n766 VDD.t1785 4.35923
R4153 VDD.n2160 VDD.n238 4.35923
R4154 VDD.n724 VDD.t3708 4.35923
R4155 VDD.n2246 VDD.t2811 4.35923
R4156 VDD.n2209 VDD.t2510 4.35923
R4157 VDD.n678 VDD.n651 4.35923
R4158 VDD.n2259 VDD.n219 4.35923
R4159 VDD.n2321 VDD.n2278 4.35923
R4160 VDD.n1474 VDD.n577 4.35914
R4161 VDD.n1505 VDD.n560 4.35914
R4162 VDD.n1557 VDD.n510 4.35914
R4163 VDD.n1529 VDD.n525 4.35914
R4164 VDD.n1597 VDD.n1596 4.35914
R4165 VDD.n1624 VDD.n1604 4.35914
R4166 VDD.n1281 VDD.n1272 4.35914
R4167 VDD.n1669 VDD.n1668 4.35914
R4168 VDD.n1718 VDD.n420 4.35914
R4169 VDD.n1689 VDD.n441 4.35914
R4170 VDD.n1775 VDD.n1774 4.35914
R4171 VDD.n1807 VDD.n1788 4.35914
R4172 VDD.n1106 VDD.n1098 4.35914
R4173 VDD.n1857 VDD.n1856 4.35914
R4174 VDD.n1900 VDD.n325 4.35914
R4175 VDD.n1949 VDD.n1948 4.35914
R4176 VDD.n1983 VDD.n1957 4.35914
R4177 VDD.n926 VDD.n919 4.35914
R4178 VDD.n2023 VDD.n2022 4.35914
R4179 VDD.n2063 VDD.n255 4.35914
R4180 VDD.n2038 VDD.n269 4.35914
R4181 VDD.n2103 VDD.n2102 4.35914
R4182 VDD.n2174 VDD.n2173 4.35914
R4183 VDD.n748 VDD.t931 4.35914
R4184 VDD.n2193 VDD.t3538 4.35914
R4185 VDD.n2228 VDD.t3943 4.35914
R4186 VDD.n2304 VDD.n2281 4.35914
R4187 VDD.n2319 VDD.n2279 4.35914
R4188 VDD.n2277 VDD.n2276 4.35914
R4189 VDD.n2261 VDD.n218 4.35914
R4190 VDD.n658 VDD.n653 4.35914
R4191 VDD.n675 VDD.n652 4.35914
R4192 VDD.n1535 VDD.t3141 4.35475
R4193 VDD.n1680 VDD.t2690 4.35475
R4194 VDD.n1495 VDD.t3432 4.35083
R4195 VDD.n1477 VDD.t3603 4.35083
R4196 VDD.n1472 VDD.t3649 4.35083
R4197 VDD.n1422 VDD.t3416 4.35083
R4198 VDD.n1572 VDD.t3284 4.35083
R4199 VDD.n1531 VDD.t3350 4.35083
R4200 VDD.n1398 VDD.t1827 4.35083
R4201 VDD.n1594 VDD.t3018 4.35083
R4202 VDD.n1623 VDD.t3543 4.35083
R4203 VDD.n1292 VDD.t3625 4.35083
R4204 VDD.n1297 VDD.t1152 4.35083
R4205 VDD.n1687 VDD.t1860 4.35083
R4206 VDD.n1806 VDD.t2953 4.35083
R4207 VDD.n1825 VDD.t3962 4.35083
R4208 VDD.n378 VDD.t4176 4.35083
R4209 VDD.n1852 VDD.t3193 4.35083
R4210 VDD.n1876 VDD.t1024 4.35083
R4211 VDD.n1934 VDD.t1518 4.35083
R4212 VDD.n1982 VDD.t993 4.35083
R4213 VDD.n1946 VDD.t4010 4.35083
R4214 VDD.n2018 VDD.t3693 4.35083
R4215 VDD.n2014 VDD.t2058 4.35083
R4216 VDD.n2055 VDD.t1623 4.35083
R4217 VDD.n2037 VDD.t1572 4.35083
R4218 VDD.n2053 VDD.t2686 4.35083
R4219 VDD.n2130 VDD.t2826 4.35083
R4220 VDD.n1290 VDD.t3619 4.34546
R4221 VDD.n1288 VDD.t974 4.34546
R4222 VDD.n1715 VDD.t2525 4.34546
R4223 VDD.n1714 VDD.t1530 4.34546
R4224 VDD.n625 VDD.t252 4.34469
R4225 VDD.n1424 VDD.t2498 4.34469
R4226 VDD.n1427 VDD.t1377 4.34469
R4227 VDD.n1437 VDD.t3058 4.34469
R4228 VDD.n1446 VDD.t1693 4.34469
R4229 VDD.n1458 VDD.t1653 4.34469
R4230 VDD.n1463 VDD.t429 4.34469
R4231 VDD.n1475 VDD.t1125 4.34469
R4232 VDD.n1481 VDD.t3908 4.34469
R4233 VDD.n1493 VDD.t2718 4.34469
R4234 VDD.n1506 VDD.t2333 4.34469
R4235 VDD.n1512 VDD.t2338 4.34469
R4236 VDD.n1509 VDD.t450 4.34469
R4237 VDD.n1521 VDD.t3412 4.34469
R4238 VDD.n1454 VDD.t4186 4.34469
R4239 VDD.n1440 VDD.t196 4.34469
R4240 VDD.n632 VDD.t869 4.34469
R4241 VDD.n1549 VDD.t3934 4.34469
R4242 VDD.n1544 VDD.t3697 4.34469
R4243 VDD.n534 VDD.t1595 4.34469
R4244 VDD.n545 VDD.t3662 4.34469
R4245 VDD.n1562 VDD.t1854 4.34469
R4246 VDD.n1404 VDD.t3286 4.34469
R4247 VDD.n1631 VDD.t793 4.34469
R4248 VDD.n1363 VDD.t3796 4.34469
R4249 VDD.n1651 VDD.t1078 4.34469
R4250 VDD.n1670 VDD.t859 4.34469
R4251 VDD.n1679 VDD.t2919 4.34469
R4252 VDD.n1795 VDD.t640 4.34469
R4253 VDD.n1840 VDD.t3067 4.34469
R4254 VDD.n1859 VDD.t64 4.34469
R4255 VDD.n1869 VDD.t1176 4.34469
R4256 VDD.n1907 VDD.t650 4.34469
R4257 VDD.n1906 VDD.t414 4.34469
R4258 VDD.n1967 VDD.t306 4.34469
R4259 VDD.n1977 VDD.t1665 4.34469
R4260 VDD.n1935 VDD.t4155 4.34469
R4261 VDD.n279 VDD.t2006 4.34469
R4262 VDD.n289 VDD.t3742 4.34469
R4263 VDD.n2168 VDD.t350 4.34469
R4264 VDD.n2175 VDD.t1009 4.34469
R4265 VDD.n2187 VDD.t4245 4.34469
R4266 VDD.n2287 VDD.t628 4.34469
R4267 VDD.n2299 VDD.t883 4.34469
R4268 VDD.n1767 VDD.t612 4.33687
R4269 VDD.n563 VDD.t2506 4.30819
R4270 VDD.n571 VDD.t903 4.30819
R4271 VDD.n584 VDD.t1408 4.30819
R4272 VDD.n606 VDD.t4019 4.30819
R4273 VDD.n1394 VDD.t3219 4.30819
R4274 VDD.n521 VDD.t865 4.30819
R4275 VDD.n503 VDD.t2785 4.30819
R4276 VDD.n484 VDD.t1929 4.30819
R4277 VDD.n1608 VDD.t2893 4.30819
R4278 VDD.n1271 VDD.t1460 4.30819
R4279 VDD.n1268 VDD.t2536 4.30819
R4280 VDD.n418 VDD.t3093 4.30819
R4281 VDD.n444 VDD.t3332 4.30819
R4282 VDD.n1793 VDD.t3000 4.30819
R4283 VDD.n383 VDD.t2122 4.30819
R4284 VDD.n1096 VDD.t2752 4.30819
R4285 VDD.n364 VDD.t2137 4.30819
R4286 VDD.n346 VDD.t3183 4.30819
R4287 VDD.n1941 VDD.t2081 4.30819
R4288 VDD.n1963 VDD.t1121 4.30819
R4289 VDD.n311 VDD.t1464 4.30819
R4290 VDD.n295 VDD.t2557 4.30819
R4291 VDD.n302 VDD.t3773 4.30819
R4292 VDD.n257 VDD.t3527 4.30819
R4293 VDD.n275 VDD.t3851 4.30819
R4294 VDD.n264 VDD.t1357 4.30819
R4295 VDD.n2111 VDD.t2435 4.30819
R4296 VDD.n1673 VDD.t1110 4.30388
R4297 VDD.n1717 VDD.t2724 4.30388
R4298 VDD.n1809 VDD.t4119 4.30388
R4299 VDD.n2138 VDD.t3124 4.30388
R4300 VDD.n1278 VDD.t1047 4.30165
R4301 VDD.n1738 VDD.t4085 4.27035
R4302 VDD.n1753 VDD.t836 4.27035
R4303 VDD.n1827 VDD.t664 4.27035
R4304 VDD.n1811 VDD.t391 4.27035
R4305 VDD.n1810 VDD.t2637 4.27035
R4306 VDD.n1766 VDD.t174 4.27035
R4307 VDD.n1107 VDD.t288 4.27035
R4308 VDD.n2101 VDD.t2283 4.27035
R4309 VDD.n2100 VDD.t1649 4.27035
R4310 VDD.n1712 VDD.t1532 4.26918
R4311 VDD.n2334 VDD.n2333 4.1315
R4312 VDD.n635 VDD.n546 4.1315
R4313 VDD.n349 VDD.t1930 3.77567
R4314 VDD.n413 VDD.t822 3.7566
R4315 VDD.n391 VDD.t148 3.7566
R4316 VDD.n382 VDD.t144 3.7566
R4317 VDD.n1779 VDD.t122 3.7566
R4318 VDD.n1780 VDD.t124 3.7566
R4319 VDD.n1091 VDD.t446 3.7566
R4320 VDD.n246 VDD.t2738 3.7566
R4321 VDD.n248 VDD.t762 3.7566
R4322 VDD.t2279 VDD.t1425 3.56594
R4323 VDD.t3349 VDD.t765 3.52369
R4324 VDD.t1709 VDD.t2384 3.47272
R4325 VDD.t729 VDD.t4059 3.47272
R4326 VDD.t4057 VDD.t4122 3.47272
R4327 VDD.t415 VDD.t1022 3.3562
R4328 VDD.n402 VDD.t1815 3.07367
R4329 VDD.n403 VDD.t1997 3.07367
R4330 VDD.n404 VDD.t1995 3.07367
R4331 VDD.n2006 VDD.n304 2.95895
R4332 VDD.n633 VDD.n612 2.85289
R4333 VDD.n1433 VDD.n604 2.85289
R4334 VDD.n1455 VDD.n590 2.85289
R4335 VDD.n1470 VDD.n579 2.85289
R4336 VDD.n1489 VDD.n569 2.85289
R4337 VDD.n1520 VDD.n550 2.85289
R4338 VDD.n1517 VDD.n553 2.85289
R4339 VDD.n1449 VDD.n594 2.85289
R4340 VDD.n628 VDD.n616 2.85289
R4341 VDD.n1548 VDD.n514 2.85289
R4342 VDD.n1542 VDD.n519 2.85289
R4343 VDD.n542 VDD.n529 2.85289
R4344 VDD.n1561 VDD.n506 2.85289
R4345 VDD.n1402 VDD.n1395 2.85289
R4346 VDD.n1362 VDD.n1342 2.85289
R4347 VDD.n1676 VDD.n461 2.85289
R4348 VDD.n1841 VDD.n376 2.85289
R4349 VDD.n1866 VDD.n363 2.85289
R4350 VDD.n1975 VDD.n1961 2.85289
R4351 VDD.n287 VDD.n273 2.85289
R4352 VDD.n2183 VDD.n233 2.85289
R4353 VDD.n2295 VDD.n2283 2.85289
R4354 VDD.n12 VDD.t221 2.8461
R4355 VDD.n25 VDD.t582 2.8461
R4356 VDD.n37 VDD.t556 2.8461
R4357 VDD.n48 VDD.t668 2.8461
R4358 VDD.n60 VDD.t264 2.8461
R4359 VDD.n72 VDD.t1758 2.8461
R4360 VDD.n84 VDD.t1312 2.8461
R4361 VDD.n96 VDD.t98 2.8461
R4362 VDD.n483 VDD.t1496 2.81423
R4363 VDD.n495 VDD.t1030 2.81423
R4364 VDD.n2105 VDD.t3126 2.81423
R4365 VDD.n1291 VDD.n1267 2.77124
R4366 VDD.n598 VDD.t1487 2.73703
R4367 VDD.n585 VDD.t3438 2.73703
R4368 VDD.n559 VDD.t2294 2.73703
R4369 VDD.n589 VDD.t2769 2.73703
R4370 VDD.n526 VDD.t1907 2.73703
R4371 VDD.n1391 VDD.t3215 2.73703
R4372 VDD.n1341 VDD.t1331 2.73703
R4373 VDD.n1610 VDD.t3835 2.73703
R4374 VDD.n481 VDD.t1102 2.73703
R4375 VDD.n491 VDD.t3122 2.73703
R4376 VDD.n493 VDD.t3027 2.73703
R4377 VDD.n497 VDD.t2439 2.73703
R4378 VDD.n1350 VDD.t3080 2.73703
R4379 VDD.n465 VDD.t3994 2.73703
R4380 VDD.n469 VDD.t1283 2.73703
R4381 VDD.n411 VDD.t3229 2.73703
R4382 VDD.n414 VDD.t2883 2.73703
R4383 VDD.n436 VDD.t2181 2.73703
R4384 VDD.n446 VDD.t2066 2.73703
R4385 VDD.n1792 VDD.t4023 2.73703
R4386 VDD.n1787 VDD.t3300 2.73703
R4387 VDD.n375 VDD.t3631 2.73703
R4388 VDD.n322 VDD.t1872 2.73703
R4389 VDD.n341 VDD.t1426 2.73703
R4390 VDD.n332 VDD.t3786 2.73703
R4391 VDD.n330 VDD.t4285 2.73703
R4392 VDD.n321 VDD.t1476 2.73703
R4393 VDD.n1958 VDD.t2377 2.73703
R4394 VDD.n316 VDD.t3500 2.73703
R4395 VDD.n297 VDD.t3601 2.73703
R4396 VDD.n270 VDD.t3981 2.73703
R4397 VDD.n2112 VDD.t3715 2.73703
R4398 VDD.n237 VDD.t2600 2.73703
R4399 VDD.n2280 VDD.t2878 2.73703
R4400 VDD.n1996 VDD.n312 2.72094
R4401 VDD.n514 VDD.t1606 2.63984
R4402 VDD.n519 VDD.t1361 2.63984
R4403 VDD.n506 VDD.t2977 2.63984
R4404 VDD.n1395 VDD.t1942 2.63984
R4405 VDD.n1342 VDD.t2263 2.63984
R4406 VDD.n376 VDD.t1296 2.63984
R4407 VDD.n512 VDD.t21 2.61116
R4408 VDD.n487 VDD.t8 2.61116
R4409 VDD.n471 VDD.t3721 2.61116
R4410 VDD.n329 VDD.t2531 2.61116
R4411 VDD.n323 VDD.t791 2.61116
R4412 VDD.n474 VDD.t801 2.55888
R4413 VDD.n477 VDD.t3730 2.55888
R4414 VDD.n478 VDD.t604 2.55888
R4415 VDD.n1274 VDD.t3728 2.55888
R4416 VDD.n2335 VDD.n213 2.55275
R4417 VDD.n133 VDD.t2352 2.44422
R4418 VDD.n132 VDD.t2022 2.44422
R4419 VDD VDD.n2336 2.41995
R4420 VDD.t2932 VDD.t1958 2.38999
R4421 VDD.n524 VDD.t2937 2.33383
R4422 VDD.n457 VDD.t3841 2.33383
R4423 VDD.n432 VDD.t1075 2.31531
R4424 VDD.n483 VDD.t3508 2.28216
R4425 VDD.n495 VDD.t2804 2.28216
R4426 VDD.n2105 VDD.t4194 2.28216
R4427 VDD.n188 VDD.n128 2.2505
R4428 VDD.n190 VDD.n189 2.2505
R4429 VDD.n191 VDD.n127 2.2505
R4430 VDD.n193 VDD.n192 2.2505
R4431 VDD.n194 VDD.n126 2.2505
R4432 VDD.n196 VDD.n195 2.2505
R4433 VDD.n197 VDD.n125 2.2505
R4434 VDD.n199 VDD.n198 2.2505
R4435 VDD.n200 VDD.n124 2.2505
R4436 VDD.n202 VDD.n201 2.2505
R4437 VDD.n203 VDD.n123 2.2505
R4438 VDD.n205 VDD.n204 2.2505
R4439 VDD.n206 VDD.n122 2.2505
R4440 VDD.n208 VDD.n207 2.2505
R4441 VDD.n209 VDD.n121 2.2505
R4442 VDD.n211 VDD.n210 2.2505
R4443 VDD.n142 VDD.t2010 2.23455
R4444 VDD.n143 VDD.t2012 2.23455
R4445 VDD.n415 VDD.t818 2.22001
R4446 VDD.n415 VDD.t820 2.22001
R4447 VDD.n389 VDD.t154 2.22001
R4448 VDD.n389 VDD.t146 2.22001
R4449 VDD.n380 VDD.t142 2.22001
R4450 VDD.n380 VDD.t152 2.22001
R4451 VDD.n1777 VDD.t118 2.22001
R4452 VDD.n1777 VDD.t42 2.22001
R4453 VDD.n1778 VDD.t120 2.22001
R4454 VDD.n1778 VDD.t622 2.22001
R4455 VDD.n402 VDD.t1819 2.22001
R4456 VDD.n403 VDD.t1821 2.22001
R4457 VDD.n404 VDD.t1823 2.22001
R4458 VDD.n1090 VDD.t816 2.22001
R4459 VDD.n1090 VDD.t824 2.22001
R4460 VDD.n249 VDD.t2735 2.22001
R4461 VDD.n249 VDD.t2736 2.22001
R4462 VDD.n250 VDD.t716 2.22001
R4463 VDD.n250 VDD.t772 2.22001
R4464 VDD.n424 VDD.t2055 2.15435
R4465 VDD.n424 VDD.t1085 2.15435
R4466 VDD.n426 VDD.t618 2.15435
R4467 VDD.n426 VDD.t808 2.15435
R4468 VDD.n428 VDD.t814 2.15435
R4469 VDD.n428 VDD.t598 2.15435
R4470 VDD.n430 VDD.t1089 2.15435
R4471 VDD.n430 VDD.t2051 2.15435
R4472 VDD.n433 VDD.t1063 2.15435
R4473 VDD.n433 VDD.t3824 2.15435
R4474 VDD.n431 VDD.t1091 2.15435
R4475 VDD.n431 VDD.t1076 2.15435
R4476 VDD.n429 VDD.t1061 2.15435
R4477 VDD.n429 VDD.t1059 2.15435
R4478 VDD.n427 VDD.t27 2.15435
R4479 VDD.n427 VDD.t1087 2.15435
R4480 VDD.n425 VDD.t1039 2.15435
R4481 VDD.n423 VDD.t38 2.15435
R4482 VDD.n423 VDD.t33 2.15435
R4483 VDD.n422 VDD.t1049 2.15435
R4484 VDD.n561 VDD.t1367 2.10455
R4485 VDD.n561 VDD.t397 2.10455
R4486 VDD.n567 VDD.t2515 2.10455
R4487 VDD.n567 VDD.t357 2.10455
R4488 VDD.n587 VDD.t4124 2.10455
R4489 VDD.n587 VDD.t1567 2.10455
R4490 VDD.n602 VDD.t1782 2.10455
R4491 VDD.n602 VDD.t4126 2.10455
R4492 VDD.n1392 VDD.t4132 2.10455
R4493 VDD.n1392 VDD.t947 2.10455
R4494 VDD.n531 VDD.t863 2.10455
R4495 VDD.n531 VDD.t393 2.10455
R4496 VDD.n518 VDD.t363 2.10455
R4497 VDD.n518 VDD.t1469 2.10455
R4498 VDD.n505 VDD.t2985 2.10455
R4499 VDD.n505 VDD.t4130 2.10455
R4500 VDD.n486 VDD.t2744 2.10455
R4501 VDD.n486 VDD.t361 2.10455
R4502 VDD.n1611 VDD.t3359 2.10455
R4503 VDD.n1611 VDD.t359 2.10455
R4504 VDD.n1273 VDD.t3025 2.10455
R4505 VDD.n1273 VDD.t4134 2.10455
R4506 VDD.n470 VDD.t395 2.10455
R4507 VDD.n470 VDD.t2357 2.10455
R4508 VDD.n1270 VDD.t3340 2.10455
R4509 VDD.n1270 VDD.t280 2.10455
R4510 VDD.n416 VDD.t4128 2.10455
R4511 VDD.n416 VDD.t3552 2.10455
R4512 VDD.n445 VDD.t1717 2.10455
R4513 VDD.n445 VDD.t399 2.10455
R4514 VDD.n1794 VDD.t3495 2.10455
R4515 VDD.n1794 VDD.t365 2.10455
R4516 VDD.n1769 VDD.t276 2.10455
R4517 VDD.n1769 VDD.t1967 2.10455
R4518 VDD.n1092 VDD.t284 2.10455
R4519 VDD.n1092 VDD.t1285 2.10455
R4520 VDD.n367 VDD.t1491 2.10455
R4521 VDD.n367 VDD.t2627 2.10455
R4522 VDD.n347 VDD.t3953 2.10455
R4523 VDD.n347 VDD.t2633 2.10455
R4524 VDD.n309 VDD.t1277 2.10455
R4525 VDD.n309 VDD.t278 2.10455
R4526 VDD.n1966 VDD.t3365 2.10455
R4527 VDD.n1966 VDD.t2631 2.10455
R4528 VDD.n314 VDD.t3476 2.10455
R4529 VDD.n314 VDD.t2619 2.10455
R4530 VDD.n296 VDD.t2190 2.10455
R4531 VDD.n296 VDD.t2617 2.10455
R4532 VDD.n305 VDD.t2621 2.10455
R4533 VDD.n305 VDD.t1507 2.10455
R4534 VDD.n254 VDD.t282 2.10455
R4535 VDD.n254 VDD.t1727 2.10455
R4536 VDD.n278 VDD.t2139 2.10455
R4537 VDD.n278 VDD.t2629 2.10455
R4538 VDD.n267 VDD.t1961 2.10455
R4539 VDD.n267 VDD.t2625 2.10455
R4540 VDD.n2113 VDD.t2034 2.10455
R4541 VDD.n2113 VDD.t2623 2.10455
R4542 VDD.n6 VDD.t227 2.0905
R4543 VDD.n19 VDD.t588 2.0905
R4544 VDD.n31 VDD.t562 2.0905
R4545 VDD.n42 VDD.t674 2.0905
R4546 VDD.n54 VDD.t270 2.0905
R4547 VDD.n66 VDD.t1744 2.0905
R4548 VDD.n78 VDD.t1318 2.0905
R4549 VDD.n90 VDD.t104 2.0905
R4550 VDD.n617 VDD.t274 2.06607
R4551 VDD.n615 VDD.t250 2.06607
R4552 VDD.n613 VDD.t244 2.06607
R4553 VDD.n612 VDD.t240 2.06607
R4554 VDD.n611 VDD.t2502 2.06607
R4555 VDD.n608 VDD.t1383 2.06607
R4556 VDD.n607 VDD.t1387 2.06607
R4557 VDD.n605 VDD.t1373 2.06607
R4558 VDD.n604 VDD.t1385 2.06607
R4559 VDD.n603 VDD.t3060 2.06607
R4560 VDD.n595 VDD.t1699 2.06607
R4561 VDD.n593 VDD.t2602 2.06607
R4562 VDD.n591 VDD.t1691 2.06607
R4563 VDD.n590 VDD.t1687 2.06607
R4564 VDD.n588 VDD.t1655 2.06607
R4565 VDD.n583 VDD.t421 2.06607
R4566 VDD.n582 VDD.t431 2.06607
R4567 VDD.n581 VDD.t425 2.06607
R4568 VDD.n579 VDD.t423 2.06607
R4569 VDD.n578 VDD.t1123 2.06607
R4570 VDD.n573 VDD.t3900 2.06607
R4571 VDD.n572 VDD.t3910 2.06607
R4572 VDD.n570 VDD.t3904 2.06607
R4573 VDD.n569 VDD.t3902 2.06607
R4574 VDD.n568 VDD.t2716 2.06607
R4575 VDD.n549 VDD.t2350 2.06607
R4576 VDD.n550 VDD.t2344 2.06607
R4577 VDD.n552 VDD.t2341 2.06607
R4578 VDD.n554 VDD.t2339 2.06607
R4579 VDD.n556 VDD.t2337 2.06607
R4580 VDD.n558 VDD.t448 2.06607
R4581 VDD.n557 VDD.t456 2.06607
R4582 VDD.n555 VDD.t452 2.06607
R4583 VDD.n553 VDD.t458 2.06607
R4584 VDD.n551 VDD.t3410 2.06607
R4585 VDD.n592 VDD.t4188 2.06607
R4586 VDD.n594 VDD.t190 2.06607
R4587 VDD.n596 VDD.t198 2.06607
R4588 VDD.n597 VDD.t192 2.06607
R4589 VDD.n599 VDD.t200 2.06607
R4590 VDD.n614 VDD.t867 2.06607
R4591 VDD.n616 VDD.t48 2.06607
R4592 VDD.n618 VDD.t52 2.06607
R4593 VDD.n619 VDD.t56 2.06607
R4594 VDD.n620 VDD.t46 2.06607
R4595 VDD.n533 VDD.t1591 2.06607
R4596 VDD.n532 VDD.t1589 2.06607
R4597 VDD.n530 VDD.t1587 2.06607
R4598 VDD.n529 VDD.t1593 2.06607
R4599 VDD.n528 VDD.t3660 2.06607
R4600 VDD.n464 VDD.t853 2.06607
R4601 VDD.n463 VDD.t572 2.06607
R4602 VDD.n462 VDD.t855 2.06607
R4603 VDD.n461 VDD.t576 2.06607
R4604 VDD.n459 VDD.t2921 2.06607
R4605 VDD.n1768 VDD.t608 2.06607
R4606 VDD.n388 VDD.t172 2.06607
R4607 VDD.n390 VDD.t178 2.06607
R4608 VDD.n392 VDD.t162 2.06607
R4609 VDD.n394 VDD.t160 2.06607
R4610 VDD.n396 VDD.t164 2.06607
R4611 VDD.n398 VDD.t166 2.06607
R4612 VDD.n399 VDD.t184 2.06607
R4613 VDD.n368 VDD.t66 2.06607
R4614 VDD.n366 VDD.t72 2.06607
R4615 VDD.n365 VDD.t86 2.06607
R4616 VDD.n363 VDD.t84 2.06607
R4617 VDD.n362 VDD.t1174 2.06607
R4618 VDD.n1965 VDD.t312 2.06607
R4619 VDD.n1964 VDD.t308 2.06607
R4620 VDD.n1962 VDD.t304 2.06607
R4621 VDD.n1961 VDD.t314 2.06607
R4622 VDD.n1960 VDD.t1669 2.06607
R4623 VDD.n277 VDD.t1874 2.06607
R4624 VDD.n276 VDD.t1919 2.06607
R4625 VDD.n274 VDD.t2004 2.06607
R4626 VDD.n273 VDD.t1876 2.06607
R4627 VDD.n272 VDD.t3738 2.06607
R4628 VDD.n236 VDD.t1015 2.06607
R4629 VDD.n235 VDD.t1011 2.06607
R4630 VDD.n234 VDD.t1007 2.06607
R4631 VDD.n233 VDD.t1017 2.06607
R4632 VDD.n232 VDD.t4249 2.06607
R4633 VDD.n2286 VDD.t658 2.06607
R4634 VDD.n2285 VDD.t654 2.06607
R4635 VDD.n2284 VDD.t626 2.06607
R4636 VDD.n2283 VDD.t630 2.06607
R4637 VDD.n2282 VDD.t887 2.06607
R4638 VDD.n512 VDD.t1393 2.03739
R4639 VDD.n487 VDD.t1275 2.03739
R4640 VDD.n471 VDD.t3255 2.03739
R4641 VDD.n329 VDD.t3678 2.03739
R4642 VDD.n323 VDD.t1051 2.03739
R4643 VDD.t2424 VDD.t2374 1.88808
R4644 VDD.n522 VDD.t799 1.84822
R4645 VDD.n522 VDD.t23 1.84822
R4646 VDD.n476 VDD.t3863 1.84822
R4647 VDD.n476 VDD.t1069 1.84822
R4648 VDD.n1666 VDD.t3392 1.84822
R4649 VDD.n1666 VDD.t29 1.84822
R4650 VDD.n474 VDD.t812 1.84822
R4651 VDD.n475 VDD.t602 1.84822
R4652 VDD.n475 VDD.t810 1.84822
R4653 VDD.n477 VDD.t3734 1.84822
R4654 VDD.n478 VDD.t610 1.84822
R4655 VDD.n1274 VDD.t1071 1.84822
R4656 VDD.n419 VDD.t3395 1.84822
R4657 VDD.n419 VDD.t31 1.84822
R4658 VDD.n417 VDD.t36 1.84822
R4659 VDD.n417 VDD.t3391 1.84822
R4660 VDD.n331 VDD.t3826 1.84822
R4661 VDD.n331 VDD.t3865 1.84822
R4662 VDD.n333 VDD.t3861 1.84822
R4663 VDD.n333 VDD.t1057 1.84822
R4664 VDD.n263 VDD.t776 1.84822
R4665 VDD.n263 VDD.t632 1.84822
R4666 VDD.n8 VDD.n5 1.80644
R4667 VDD.n9 VDD.n4 1.80644
R4668 VDD.n10 VDD.n3 1.80644
R4669 VDD.n11 VDD.n2 1.80644
R4670 VDD.n21 VDD.n18 1.80644
R4671 VDD.n22 VDD.n17 1.80644
R4672 VDD.n23 VDD.n16 1.80644
R4673 VDD.n24 VDD.n15 1.80644
R4674 VDD.n33 VDD.n30 1.80644
R4675 VDD.n34 VDD.n29 1.80644
R4676 VDD.n35 VDD.n28 1.80644
R4677 VDD.n36 VDD.n27 1.80644
R4678 VDD.n44 VDD.n41 1.80644
R4679 VDD.n45 VDD.n40 1.80644
R4680 VDD.n46 VDD.n39 1.80644
R4681 VDD.n47 VDD.n38 1.80644
R4682 VDD.n56 VDD.n53 1.80644
R4683 VDD.n57 VDD.n52 1.80644
R4684 VDD.n58 VDD.n51 1.80644
R4685 VDD.n59 VDD.n50 1.80644
R4686 VDD.n68 VDD.n65 1.80644
R4687 VDD.n69 VDD.n64 1.80644
R4688 VDD.n70 VDD.n63 1.80644
R4689 VDD.n71 VDD.n62 1.80644
R4690 VDD.n80 VDD.n77 1.80644
R4691 VDD.n81 VDD.n76 1.80644
R4692 VDD.n82 VDD.n75 1.80644
R4693 VDD.n83 VDD.n74 1.80644
R4694 VDD.n92 VDD.n89 1.80644
R4695 VDD.n93 VDD.n88 1.80644
R4696 VDD.n94 VDD.n87 1.80644
R4697 VDD.n95 VDD.n86 1.80644
R4698 VDD.n575 VDD.t3403 1.75837
R4699 VDD.n547 VDD.t3629 1.75837
R4700 VDD.n496 VDD.t1238 1.75837
R4701 VDD.n1348 VDD.t930 1.75837
R4702 VDD.n1347 VDD.t1661 1.75837
R4703 VDD.n360 VDD.t1258 1.75837
R4704 VDD.n317 VDD.t2475 1.75837
R4705 VDD.n313 VDD.t1964 1.75837
R4706 VDD.n917 VDD.t3330 1.75837
R4707 VDD.n2110 VDD.t1677 1.75837
R4708 VDD.n598 VDD.t1944 1.73383
R4709 VDD.n585 VDD.t1602 1.73383
R4710 VDD.n559 VDD.t3769 1.73383
R4711 VDD.n589 VDD.t2975 1.73383
R4712 VDD.n526 VDD.t62 1.73383
R4713 VDD.n1391 VDD.t1704 1.73383
R4714 VDD.n1341 VDD.t2765 1.73383
R4715 VDD.n1610 VDD.t1108 1.73383
R4716 VDD.n481 VDD.t1514 1.73383
R4717 VDD.n491 VDD.t3607 1.73383
R4718 VDD.n493 VDD.t1509 1.73383
R4719 VDD.n497 VDD.t4166 1.73383
R4720 VDD.n1350 VDD.t2411 1.73383
R4721 VDD.n465 VDD.t1264 1.73383
R4722 VDD.n469 VDD.t3777 1.73383
R4723 VDD.n411 VDD.t336 1.73383
R4724 VDD.n414 VDD.t1167 1.73383
R4725 VDD.n436 VDD.t3245 1.73383
R4726 VDD.n446 VDD.t2605 1.73383
R4727 VDD.n1792 VDD.t3243 1.73383
R4728 VDD.n1787 VDD.t1223 1.73383
R4729 VDD.n375 VDD.t917 1.73383
R4730 VDD.n322 VDD.t1775 1.73383
R4731 VDD.n341 VDD.t2280 1.73383
R4732 VDD.n332 VDD.t4210 1.73383
R4733 VDD.n330 VDD.t2596 1.73383
R4734 VDD.n321 VDD.t1797 1.73383
R4735 VDD.n1958 VDD.t1288 1.73383
R4736 VDD.n316 VDD.t1466 1.73383
R4737 VDD.n297 VDD.t2077 1.73383
R4738 VDD.n270 VDD.t1262 1.73383
R4739 VDD.n2112 VDD.t2427 1.73383
R4740 VDD.n237 VDD.t2100 1.73383
R4741 VDD.n2280 VDD.t3702 1.73383
R4742 VDD.n312 VDD.t1204 1.72898
R4743 VDD.n2334 VDD.n214 1.7051
R4744 VDD.n636 VDD.n635 1.7051
R4745 VDD.n413 VDD.t4095 1.67844
R4746 VDD.n391 VDD.t842 1.67844
R4747 VDD.n382 VDD.t690 1.67844
R4748 VDD.n1779 VDD.t353 1.67844
R4749 VDD.n1780 VDD.t2609 1.67844
R4750 VDD.n1091 VDD.t290 1.67844
R4751 VDD.n246 VDD.t2289 1.67844
R4752 VDD.n248 VDD.t1645 1.67844
R4753 VDD.n99 VDD.n98 1.52602
R4754 VDD.n400 VDD.t186 1.52029
R4755 VDD.n1267 VDD.t3621 1.49844
R4756 VDD.n1267 VDD.t3623 1.49844
R4757 VDD.n460 VDD.t2407 1.49844
R4758 VDD.n460 VDD.t3820 1.49844
R4759 VDD.n472 VDD.t3235 1.49844
R4760 VDD.n472 VDD.t3926 1.49844
R4761 VDD.n434 VDD.t3818 1.49844
R4762 VDD.n434 VDD.t3022 1.49844
R4763 VDD.n443 VDD.t926 1.49844
R4764 VDD.n443 VDD.t3105 1.49844
R4765 VDD.n335 VDD.t3497 1.49844
R4766 VDD.n335 VDD.t2096 1.49844
R4767 VDD.n1951 VDD.t2312 1.49844
R4768 VDD.n1951 VDD.t2563 1.49844
R4769 VDD.n1956 VDD.t964 1.49844
R4770 VDD.n1956 VDD.t3816 1.49844
R4771 VDD.n306 VDD.t2413 1.49844
R4772 VDD.n306 VDD.t3723 1.49844
R4773 VDD.n298 VDD.t3213 1.49844
R4774 VDD.n298 VDD.t3107 1.49844
R4775 VDD.n260 VDD.t3651 1.49844
R4776 VDD.n260 VDD.t3151 1.49844
R4777 VDD.n617 VDD.t246 1.4923
R4778 VDD.n615 VDD.t242 1.4923
R4779 VDD.n613 VDD.t248 1.4923
R4780 VDD.n612 VDD.t2496 1.4923
R4781 VDD.n611 VDD.t2500 1.4923
R4782 VDD.n608 VDD.t1375 1.4923
R4783 VDD.n607 VDD.t1381 1.4923
R4784 VDD.n605 VDD.t1379 1.4923
R4785 VDD.n604 VDD.t3062 1.4923
R4786 VDD.n603 VDD.t3063 1.4923
R4787 VDD.n595 VDD.t1689 1.4923
R4788 VDD.n593 VDD.t1697 1.4923
R4789 VDD.n591 VDD.t1695 1.4923
R4790 VDD.n590 VDD.t1657 1.4923
R4791 VDD.n588 VDD.t1659 1.4923
R4792 VDD.n583 VDD.t427 1.4923
R4793 VDD.n582 VDD.t435 1.4923
R4794 VDD.n581 VDD.t433 1.4923
R4795 VDD.n579 VDD.t1127 1.4923
R4796 VDD.n578 VDD.t1129 1.4923
R4797 VDD.n573 VDD.t3906 1.4923
R4798 VDD.n572 VDD.t3898 1.4923
R4799 VDD.n570 VDD.t3896 1.4923
R4800 VDD.n569 VDD.t2712 1.4923
R4801 VDD.n568 VDD.t2714 1.4923
R4802 VDD.n549 VDD.t2335 1.4923
R4803 VDD.n550 VDD.t2348 1.4923
R4804 VDD.n552 VDD.t2346 1.4923
R4805 VDD.n554 VDD.t2342 1.4923
R4806 VDD.n556 VDD.t2336 1.4923
R4807 VDD.n558 VDD.t620 1.4923
R4808 VDD.n557 VDD.t454 1.4923
R4809 VDD.n555 VDD.t460 1.4923
R4810 VDD.n553 VDD.t3411 1.4923
R4811 VDD.n551 VDD.t3409 1.4923
R4812 VDD.n592 VDD.t4192 1.4923
R4813 VDD.n594 VDD.t4190 1.4923
R4814 VDD.n596 VDD.t202 1.4923
R4815 VDD.n597 VDD.t194 1.4923
R4816 VDD.n599 VDD.t204 1.4923
R4817 VDD.n614 VDD.t873 1.4923
R4818 VDD.n616 VDD.t871 1.4923
R4819 VDD.n618 VDD.t60 1.4923
R4820 VDD.n619 VDD.t50 1.4923
R4821 VDD.n620 VDD.t54 1.4923
R4822 VDD.n514 VDD.t3932 1.4923
R4823 VDD.n516 VDD.t1363 1.4923
R4824 VDD.n516 VDD.t3029 1.4923
R4825 VDD.n519 VDD.t3695 1.4923
R4826 VDD.n520 VDD.t692 1.4923
R4827 VDD.n520 VDD.t18 1.4923
R4828 VDD.n533 VDD.t1596 1.4923
R4829 VDD.n532 VDD.t1598 1.4923
R4830 VDD.n530 VDD.t1600 1.4923
R4831 VDD.n529 VDD.t3664 1.4923
R4832 VDD.n528 VDD.t3658 1.4923
R4833 VDD.n509 VDD.t3802 1.4923
R4834 VDD.n509 VDD.t3032 1.4923
R4835 VDD.n506 VDD.t1856 1.4923
R4836 VDD.n1396 VDD.t2672 1.4923
R4837 VDD.n1396 VDD.t2224 1.4923
R4838 VDD.n1395 VDD.t3288 1.4923
R4839 VDD.n1344 VDD.t1940 1.4923
R4840 VDD.n1344 VDD.t2227 1.4923
R4841 VDD.n1342 VDD.t3798 1.4923
R4842 VDD.n464 VDD.t851 1.4923
R4843 VDD.n463 VDD.t574 1.4923
R4844 VDD.n462 VDD.t857 1.4923
R4845 VDD.n461 VDD.t2915 1.4923
R4846 VDD.n459 VDD.t2917 1.4923
R4847 VDD.n412 VDD.t4087 1.4923
R4848 VDD.n412 VDD.t4091 1.4923
R4849 VDD.n410 VDD.t4083 1.4923
R4850 VDD.n410 VDD.t4093 1.4923
R4851 VDD.n408 VDD.t4089 1.4923
R4852 VDD.n408 VDD.t4081 1.4923
R4853 VDD.n397 VDD.t830 1.4923
R4854 VDD.n397 VDD.t840 1.4923
R4855 VDD.n395 VDD.t828 1.4923
R4856 VDD.n395 VDD.t834 1.4923
R4857 VDD.n393 VDD.t838 1.4923
R4858 VDD.n393 VDD.t832 1.4923
R4859 VDD.n1768 VDD.t600 1.4923
R4860 VDD.n384 VDD.t700 1.4923
R4861 VDD.n384 VDD.t688 1.4923
R4862 VDD.n385 VDD.t698 1.4923
R4863 VDD.n385 VDD.t662 1.4923
R4864 VDD.n386 VDD.t696 1.4923
R4865 VDD.n386 VDD.t660 1.4923
R4866 VDD.n1781 VDD.t320 1.4923
R4867 VDD.n1781 VDD.t389 1.4923
R4868 VDD.n1783 VDD.t355 1.4923
R4869 VDD.n1783 VDD.t387 1.4923
R4870 VDD.n1785 VDD.t348 1.4923
R4871 VDD.n1785 VDD.t322 1.4923
R4872 VDD.n1786 VDD.t2639 1.4923
R4873 VDD.n1786 VDD.t2613 1.4923
R4874 VDD.n1784 VDD.t2607 1.4923
R4875 VDD.n1784 VDD.t2615 1.4923
R4876 VDD.n1782 VDD.t2611 1.4923
R4877 VDD.n1782 VDD.t2635 1.4923
R4878 VDD.n388 VDD.t176 1.4923
R4879 VDD.n390 VDD.t188 1.4923
R4880 VDD.n392 VDD.t158 1.4923
R4881 VDD.n394 VDD.t168 1.4923
R4882 VDD.n396 VDD.t170 1.4923
R4883 VDD.n398 VDD.t180 1.4923
R4884 VDD.n399 VDD.t182 1.4923
R4885 VDD.n376 VDD.t3065 1.4923
R4886 VDD.n374 VDD.t1221 1.4923
R4887 VDD.n374 VDD.t1034 1.4923
R4888 VDD.n368 VDD.t417 1.4923
R4889 VDD.n366 VDD.t70 1.4923
R4890 VDD.n365 VDD.t68 1.4923
R4891 VDD.n363 VDD.t1172 1.4923
R4892 VDD.n362 VDD.t1178 1.4923
R4893 VDD.n1095 VDD.t296 1.4923
R4894 VDD.n1095 VDD.t300 1.4923
R4895 VDD.n1094 VDD.t294 1.4923
R4896 VDD.n1094 VDD.t286 1.4923
R4897 VDD.n1093 VDD.t298 1.4923
R4898 VDD.n1093 VDD.t292 1.4923
R4899 VDD.n1965 VDD.t316 1.4923
R4900 VDD.n1964 VDD.t302 1.4923
R4901 VDD.n1962 VDD.t310 1.4923
R4902 VDD.n1961 VDD.t1667 1.4923
R4903 VDD.n1960 VDD.t1671 1.4923
R4904 VDD.n277 VDD.t1878 1.4923
R4905 VDD.n276 VDD.t2002 1.4923
R4906 VDD.n274 VDD.t1921 1.4923
R4907 VDD.n273 VDD.t3740 1.4923
R4908 VDD.n272 VDD.t3744 1.4923
R4909 VDD.n2099 VDD.t2286 1.4923
R4910 VDD.n2099 VDD.t2287 1.4923
R4911 VDD.n242 VDD.t1647 1.4923
R4912 VDD.n242 VDD.t1639 1.4923
R4913 VDD.n241 VDD.t2284 1.4923
R4914 VDD.n241 VDD.t2290 1.4923
R4915 VDD.n245 VDD.t1651 1.4923
R4916 VDD.n245 VDD.t1643 1.4923
R4917 VDD.n244 VDD.t2288 1.4923
R4918 VDD.n244 VDD.t2281 1.4923
R4919 VDD.n247 VDD.t1637 1.4923
R4920 VDD.n247 VDD.t1641 1.4923
R4921 VDD.n236 VDD.t1019 1.4923
R4922 VDD.n235 VDD.t1005 1.4923
R4923 VDD.n234 VDD.t1013 1.4923
R4924 VDD.n233 VDD.t4247 1.4923
R4925 VDD.n232 VDD.t4243 1.4923
R4926 VDD.n2286 VDD.t666 1.4923
R4927 VDD.n2285 VDD.t624 1.4923
R4928 VDD.n2284 VDD.t656 1.4923
R4929 VDD.n2283 VDD.t885 1.4923
R4930 VDD.n2282 VDD.t889 1.4923
R4931 VDD.n2127 VDD.n2109 1.44746
R4932 VDD.n304 VDD.t3754 1.43493
R4933 VDD.n565 VDD.t745 1.39717
R4934 VDD.n574 VDD.t768 1.39717
R4935 VDD.n580 VDD.t770 1.39717
R4936 VDD.n609 VDD.t737 1.39717
R4937 VDD.n1397 VDD.t740 1.39717
R4938 VDD.n523 VDD.t742 1.39717
R4939 VDD.n501 VDD.t705 1.39717
R4940 VDD.n1590 VDD.t510 1.39717
R4941 VDD.n1606 VDD.t516 1.39717
R4942 VDD.n1266 VDD.t760 1.39717
R4943 VDD.n442 VDD.t464 1.39717
R4944 VDD.n1790 VDD.t521 1.39717
R4945 VDD.n387 VDD.t524 1.39717
R4946 VDD.n1100 VDD.t728 1.39717
R4947 VDD.n1854 VDD.t500 1.39717
R4948 VDD.n344 VDD.t514 1.39717
R4949 VDD.n315 VDD.t730 1.39717
R4950 VDD.n1959 VDD.t502 1.39717
R4951 VDD.n1942 VDD.t540 1.39717
R4952 VDD.n292 VDD.t487 1.39717
R4953 VDD.n300 VDD.t495 1.39717
R4954 VDD.n259 VDD.t512 1.39717
R4955 VDD.n271 VDD.t470 1.39717
R4956 VDD.n261 VDD.t526 1.39717
R4957 VDD.n2108 VDD.t489 1.39717
R4958 VDD.n1269 VDD.t712 1.34263
R4959 VDD.n421 VDD.t707 1.34263
R4960 VDD.n1877 VDD.n342 1.32014
R4961 VDD.n1482 VDD.n546 1.31506
R4962 VDD.n2333 VDD.n2332 1.31506
R4963 VDD.n636 VDD.n499 1.31506
R4964 VDD.n2254 VDD.n214 1.31506
R4965 VDD.t513 VDD.t2279 1.04916
R4966 VDD.n213 VDD.n212 0.976933
R4967 VDD.n49 VDD.n37 0.928233
R4968 VDD.n2336 VDD.n2335 0.8455
R4969 VDD.n1409 VDD.n1408 0.8405
R4970 VDD.t996 VDD.n349 0.839426
R4971 VDD.t786 VDD.t2424 0.839426
R4972 VDD.n109 VDD.n108 0.808608
R4973 VDD.n61 VDD.n49 0.803758
R4974 VDD.n73 VDD.n61 0.803758
R4975 VDD.n85 VDD.n73 0.803758
R4976 VDD.n97 VDD.n85 0.803758
R4977 VDD.n1990 VDD.n1989 0.788
R4978 VDD.n1499 VDD.n1498 0.78425
R4979 VDD.n1305 VDD.n1304 0.7625
R4980 VDD.n1988 VDD.n1987 0.761
R4981 VDD.n1694 VDD.n1693 0.743
R4982 VDD.n1632 VDD.n1631 0.72275
R4983 VDD.n1882 VDD.n1881 0.69275
R4984 VDD.n1692 VDD.n1691 0.68225
R4985 VDD.n1880 VDD.n1879 0.67775
R4986 VDD.n115 VDD.t367 0.6505
R4987 VDD.n115 VDD.t371 0.6505
R4988 VDD.n114 VDD.t369 0.6505
R4989 VDD.n114 VDD.t383 0.6505
R4990 VDD.n110 VDD.t381 0.6505
R4991 VDD.n110 VDD.t385 0.6505
R4992 VDD.n111 VDD.t375 0.6505
R4993 VDD.n111 VDD.t379 0.6505
R4994 VDD.n182 VDD.t334 0.6505
R4995 VDD.n182 VDD.t330 0.6505
R4996 VDD.n181 VDD.t326 0.6505
R4997 VDD.n181 VDD.t328 0.6505
R4998 VDD.n176 VDD.t344 0.6505
R4999 VDD.n176 VDD.t346 0.6505
R5000 VDD.n177 VDD.t342 0.6505
R5001 VDD.n177 VDD.t338 0.6505
R5002 VDD.n5 VDD.t223 0.6505
R5003 VDD.n5 VDD.t235 0.6505
R5004 VDD.n4 VDD.t217 0.6505
R5005 VDD.n4 VDD.t229 0.6505
R5006 VDD.n3 VDD.t219 0.6505
R5007 VDD.n3 VDD.t231 0.6505
R5008 VDD.n2 VDD.t233 0.6505
R5009 VDD.n2 VDD.t225 0.6505
R5010 VDD.n18 VDD.t584 0.6505
R5011 VDD.n18 VDD.t596 0.6505
R5012 VDD.n17 VDD.t578 0.6505
R5013 VDD.n17 VDD.t590 0.6505
R5014 VDD.n16 VDD.t580 0.6505
R5015 VDD.n16 VDD.t592 0.6505
R5016 VDD.n15 VDD.t594 0.6505
R5017 VDD.n15 VDD.t586 0.6505
R5018 VDD.n30 VDD.t570 0.6505
R5019 VDD.n30 VDD.t558 0.6505
R5020 VDD.n29 VDD.t554 0.6505
R5021 VDD.n29 VDD.t564 0.6505
R5022 VDD.n28 VDD.t560 0.6505
R5023 VDD.n28 VDD.t566 0.6505
R5024 VDD.n27 VDD.t568 0.6505
R5025 VDD.n27 VDD.t552 0.6505
R5026 VDD.n41 VDD.t682 0.6505
R5027 VDD.n41 VDD.t670 0.6505
R5028 VDD.n40 VDD.t686 0.6505
R5029 VDD.n40 VDD.t676 0.6505
R5030 VDD.n39 VDD.t672 0.6505
R5031 VDD.n39 VDD.t678 0.6505
R5032 VDD.n38 VDD.t680 0.6505
R5033 VDD.n38 VDD.t684 0.6505
R5034 VDD.n53 VDD.t258 0.6505
R5035 VDD.n53 VDD.t266 0.6505
R5036 VDD.n52 VDD.t262 0.6505
R5037 VDD.n52 VDD.t272 0.6505
R5038 VDD.n51 VDD.t268 0.6505
R5039 VDD.n51 VDD.t254 0.6505
R5040 VDD.n50 VDD.t256 0.6505
R5041 VDD.n50 VDD.t260 0.6505
R5042 VDD.n65 VDD.t1760 0.6505
R5043 VDD.n65 VDD.t1752 0.6505
R5044 VDD.n64 VDD.t1754 0.6505
R5045 VDD.n64 VDD.t1746 0.6505
R5046 VDD.n63 VDD.t1756 0.6505
R5047 VDD.n63 VDD.t1748 0.6505
R5048 VDD.n62 VDD.t1750 0.6505
R5049 VDD.n62 VDD.t1742 0.6505
R5050 VDD.n77 VDD.t1314 0.6505
R5051 VDD.n77 VDD.t1306 0.6505
R5052 VDD.n76 VDD.t1308 0.6505
R5053 VDD.n76 VDD.t1320 0.6505
R5054 VDD.n75 VDD.t1310 0.6505
R5055 VDD.n75 VDD.t1302 0.6505
R5056 VDD.n74 VDD.t1304 0.6505
R5057 VDD.n74 VDD.t1316 0.6505
R5058 VDD.n89 VDD.t100 0.6505
R5059 VDD.n89 VDD.t92 0.6505
R5060 VDD.n88 VDD.t94 0.6505
R5061 VDD.n88 VDD.t106 0.6505
R5062 VDD.n87 VDD.t96 0.6505
R5063 VDD.n87 VDD.t88 0.6505
R5064 VDD.n86 VDD.t90 0.6505
R5065 VDD.n86 VDD.t102 0.6505
R5066 VDD.n1180 VDD.n1179 0.64625
R5067 VDD.n1502 VDD.n1501 0.6455
R5068 VDD.n1566 VDD.n1565 0.6455
R5069 VDD.n1798 VDD.n1797 0.6455
R5070 VDD.n2028 VDD.n2027 0.6455
R5071 VDD.n1852 VDD.n1851 0.635
R5072 VDD.n134 VDD.n133 0.635
R5073 VDD.n2045 VDD.n2044 0.629
R5074 VDD.n2031 VDD.n2030 0.62225
R5075 VDD.n1886 VDD.n1885 0.6185
R5076 VDD.n1585 VDD.n1584 0.61625
R5077 VDD.n1541 VDD.n1540 0.6155
R5078 VDD.n1630 VDD.n1629 0.5885
R5079 VDD.n1546 VDD.n1545 0.5825
R5080 VDD.n98 VDD.n97 0.574192
R5081 VDD.n1286 VDD.n1285 0.56525
R5082 VDD.n1412 VDD.n1411 0.55625
R5083 VDD.n2122 VDD.n2121 0.5555
R5084 VDD.n1996 VDD.n1995 0.5375
R5085 VDD.n1414 VDD.n1413 0.53075
R5086 VDD.n1104 VDD.n1103 0.53075
R5087 VDD.n1848 VDD.n1847 0.53075
R5088 VDD.n1843 VDD.n1842 0.5285
R5089 VDD.n929 VDD.n928 0.527
R5090 VDD.n355 VDD.n354 0.518
R5091 VDD.n1356 VDD.n1355 0.5105
R5092 VDD.n1547 VDD.n1546 0.50825
R5093 VDD.n1615 VDD.n1614 0.506
R5094 VDD.n2005 VDD.n2004 0.5045
R5095 VDD.n1900 VDD.n1899 0.50075
R5096 VDD.n2018 VDD.n2017 0.50075
R5097 VDD.n1560 VDD.n1559 0.497
R5098 VDD.n450 VDD.n449 0.497
R5099 VDD.n1939 VDD.n1938 0.497
R5100 VDD.n2135 VDD.n2134 0.497
R5101 VDD.n2011 VDD.n2010 0.49025
R5102 VDD.n1665 VDD.n1664 0.4865
R5103 VDD.n134 VDD.n132 0.4865
R5104 VDD.n1579 VDD.n1578 0.479
R5105 VDD.n1583 VDD.n1582 0.47225
R5106 VDD.n1986 VDD.n1985 0.4655
R5107 VDD.n1802 VDD.n1801 0.4625
R5108 VDD.n358 VDD.n357 0.4625
R5109 VDD.n1400 VDD.n1399 0.45425
R5110 VDD.n1696 VDD.n1695 0.44975
R5111 VDD.n1619 VDD.n1618 0.44375
R5112 VDD.n1419 VDD.n1418 0.4415
R5113 VDD.n1418 VDD.n1372 0.4415
R5114 VDD.n1372 VDD.n1332 0.4415
R5115 VDD.n1332 VDD.n1247 0.4415
R5116 VDD.n1247 VDD.n1206 0.4415
R5117 VDD.n1206 VDD.n1160 0.4415
R5118 VDD.n1160 VDD.n1074 0.4415
R5119 VDD.n1074 VDD.n1027 0.4415
R5120 VDD.n1027 VDD.n980 0.4415
R5121 VDD.n980 VDD.n900 0.4415
R5122 VDD.n900 VDD.n853 0.4415
R5123 VDD.n853 VDD.n806 0.4415
R5124 VDD.n806 VDD.n727 0.4415
R5125 VDD.n727 VDD.n680 0.4415
R5126 VDD.n1525 VDD.n1524 0.4415
R5127 VDD.n1525 VDD.n456 0.4415
R5128 VDD.n1683 VDD.n456 0.4415
R5129 VDD.n1684 VDD.n1683 0.4415
R5130 VDD.n1684 VDD.n359 0.4415
R5131 VDD.n1871 VDD.n359 0.4415
R5132 VDD.n1872 VDD.n1871 0.4415
R5133 VDD.n1872 VDD.n291 0.4415
R5134 VDD.n2032 VDD.n291 0.4415
R5135 VDD.n2033 VDD.n2032 0.4415
R5136 VDD.n2033 VDD.n230 0.4415
R5137 VDD.n2189 VDD.n230 0.4415
R5138 VDD.n2190 VDD.n2189 0.4415
R5139 VDD.n2190 VDD.n215 0.4415
R5140 VDD.n1482 VDD.n480 0.4415
R5141 VDD.n1642 VDD.n480 0.4415
R5142 VDD.n1643 VDD.n1642 0.4415
R5143 VDD.n1643 VDD.n379 0.4415
R5144 VDD.n1836 VDD.n379 0.4415
R5145 VDD.n1837 VDD.n1836 0.4415
R5146 VDD.n1837 VDD.n308 0.4415
R5147 VDD.n2000 VDD.n308 0.4415
R5148 VDD.n2001 VDD.n2000 0.4415
R5149 VDD.n2001 VDD.n240 0.4415
R5150 VDD.n2150 VDD.n240 0.4415
R5151 VDD.n2151 VDD.n2150 0.4415
R5152 VDD.n2151 VDD.n216 0.4415
R5153 VDD.n2332 VDD.n216 0.4415
R5154 VDD.n1575 VDD.n499 0.4415
R5155 VDD.n1576 VDD.n1575 0.4415
R5156 VDD.n1576 VDD.n406 0.4415
R5157 VDD.n1741 VDD.n406 0.4415
R5158 VDD.n1742 VDD.n1741 0.4415
R5159 VDD.n1742 VDD.n319 0.4415
R5160 VDD.n1920 VDD.n319 0.4415
R5161 VDD.n1921 VDD.n1920 0.4415
R5162 VDD.n1921 VDD.n252 0.4415
R5163 VDD.n2081 VDD.n252 0.4415
R5164 VDD.n2082 VDD.n2081 0.4415
R5165 VDD.n2082 VDD.n221 0.4415
R5166 VDD.n2253 VDD.n221 0.4415
R5167 VDD.n2254 VDD.n2253 0.4415
R5168 VDD.n2055 VDD.n2054 0.4355
R5169 VDD.n1587 VDD.n1586 0.43325
R5170 VDD.n1898 VDD.n1897 0.43325
R5171 VDD.n1361 VDD.n1360 0.43025
R5172 VDD.n2004 VDD.n2003 0.42575
R5173 VDD.n1849 VDD.n1848 0.422
R5174 VDD.n1851 VDD.n1850 0.422
R5175 VDD.n1905 VDD.n1904 0.4205
R5176 VDD.n1357 VDD.n1356 0.4175
R5177 VDD.n924 VDD.n923 0.41525
R5178 VDD.n1558 VDD.n1557 0.4145
R5179 VDD.n1578 VDD.n1577 0.413
R5180 VDD.n1591 VDD.n482 0.4115
R5181 VDD.n1661 VDD.n1660 0.41075
R5182 VDD.n2060 VDD.n2059 0.41075
R5183 VDD.n1653 VDD.n1652 0.4025
R5184 VDD.n1354 VDD.n1353 0.39425
R5185 VDD.n1663 VDD.n1662 0.3905
R5186 VDD.n1582 VDD.n1581 0.3845
R5187 VDD.n2016 VDD.n2015 0.3815
R5188 VDD.n2128 VDD.n2127 0.37625
R5189 VDD.n1637 VDD.n1636 0.3755
R5190 VDD.n1846 VDD.n1845 0.3725
R5191 VDD.n2009 VDD.n2008 0.3725
R5192 VDD.n1353 VDD.n1352 0.36875
R5193 VDD.n1529 VDD.n1528 0.3665
R5194 VDD.n1884 VDD.n1883 0.36575
R5195 VDD.n1628 VDD.n1627 0.36275
R5196 VDD.n2025 VDD.n2024 0.3605
R5197 VDD.n212 VDD.n211 0.35997
R5198 VDD.n188 VDD.n187 0.359916
R5199 VDD.n1835 VDD.n381 0.356
R5200 VDD.n1463 VDD.n1462 0.3515
R5201 VDD.n2137 VDD.n2136 0.35075
R5202 VDD.n925 VDD.n924 0.34775
R5203 VDD.n1985 VDD.n1984 0.34175
R5204 VDD.n2166 VDD.n2165 0.34175
R5205 VDD.n1618 VDD.n1617 0.341
R5206 VDD.n1850 VDD.n1849 0.341
R5207 VDD.n2102 VDD.n2101 0.3395
R5208 VDD.n2127 VDD.n2126 0.3395
R5209 VDD.n1912 VDD.n1911 0.33725
R5210 VDD.n1930 VDD.n1929 0.33725
R5211 VDD.n1428 VDD.n1427 0.3365
R5212 VDD.n1433 VDD.n1432 0.3365
R5213 VDD.n1468 VDD.n1467 0.3365
R5214 VDD.n1489 VDD.n1488 0.3365
R5215 VDD.n1385 VDD.n1384 0.3365
R5216 VDD.n1382 VDD.n1381 0.3365
R5217 VDD.n1379 VDD.n1378 0.3365
R5218 VDD.n543 VDD.n542 0.3365
R5219 VDD.n1339 VDD.n1338 0.3365
R5220 VDD.n1338 VDD.n1337 0.3365
R5221 VDD.n1337 VDD.n1336 0.3365
R5222 VDD.n1336 VDD.n1335 0.3365
R5223 VDD.n1335 VDD.n1334 0.3365
R5224 VDD.n1334 VDD.n1333 0.3365
R5225 VDD.n1368 VDD.n1367 0.3365
R5226 VDD.n1365 VDD.n1364 0.3365
R5227 VDD.n1676 VDD.n1675 0.3365
R5228 VDD.n1675 VDD.n1674 0.3365
R5229 VDD.n1225 VDD.n1224 0.3365
R5230 VDD.n1224 VDD.n1223 0.3365
R5231 VDD.n1223 VDD.n1222 0.3365
R5232 VDD.n1222 VDD.n1221 0.3365
R5233 VDD.n1221 VDD.n407 0.3365
R5234 VDD.n1732 VDD.n1731 0.3365
R5235 VDD.n1182 VDD.n1181 0.3365
R5236 VDD.n1830 VDD.n1829 0.3365
R5237 VDD.n1120 VDD.n1119 0.3365
R5238 VDD.n1119 VDD.n1118 0.3365
R5239 VDD.n1118 VDD.n1117 0.3365
R5240 VDD.n1110 VDD.n1109 0.3365
R5241 VDD.n1860 VDD.n1859 0.3365
R5242 VDD.n1976 VDD.n1975 0.3365
R5243 VDD.n932 VDD.n931 0.3365
R5244 VDD.n931 VDD.n930 0.3365
R5245 VDD.n2073 VDD.n2072 0.3365
R5246 VDD.n2072 VDD.n2071 0.3365
R5247 VDD.n2071 VDD.n2070 0.3365
R5248 VDD.n2070 VDD.n2069 0.3365
R5249 VDD.n2069 VDD.n2068 0.3365
R5250 VDD.n2068 VDD.n2067 0.3365
R5251 VDD.n2042 VDD.n2041 0.3365
R5252 VDD.n288 VDD.n287 0.3365
R5253 VDD.n2091 VDD.n2090 0.3365
R5254 VDD.n2092 VDD.n2091 0.3365
R5255 VDD.n2093 VDD.n2092 0.3365
R5256 VDD.n2094 VDD.n2093 0.3365
R5257 VDD.n2095 VDD.n2094 0.3365
R5258 VDD.n2096 VDD.n2095 0.3365
R5259 VDD.n2097 VDD.n2096 0.3365
R5260 VDD.n2098 VDD.n2097 0.3365
R5261 VDD.n2101 VDD.n2100 0.3365
R5262 VDD.n2100 VDD.n243 0.3365
R5263 VDD.n2148 VDD.n2147 0.3365
R5264 VDD.n2147 VDD.n2146 0.3365
R5265 VDD.n2145 VDD.n2144 0.3365
R5266 VDD.n2118 VDD.n2117 0.3365
R5267 VDD.n2117 VDD.n2116 0.3365
R5268 VDD.n2158 VDD.n2157 0.3365
R5269 VDD.n2159 VDD.n2158 0.3365
R5270 VDD.n2164 VDD.n2163 0.3365
R5271 VDD.n2172 VDD.n231 0.3365
R5272 VDD.n2200 VDD.n2199 0.3365
R5273 VDD.n229 VDD.n228 0.3365
R5274 VDD.n228 VDD.n227 0.3365
R5275 VDD.n227 VDD.n226 0.3365
R5276 VDD.n226 VDD.n225 0.3365
R5277 VDD.n225 VDD.n224 0.3365
R5278 VDD.n224 VDD.n223 0.3365
R5279 VDD.n677 VDD.n676 0.3365
R5280 VDD.n657 VDD.n656 0.3365
R5281 VDD.n656 VDD.n655 0.3365
R5282 VDD.n655 VDD.n654 0.3365
R5283 VDD.n654 VDD.n220 0.3365
R5284 VDD.n2257 VDD.n2256 0.3365
R5285 VDD.n2258 VDD.n2257 0.3365
R5286 VDD.n2263 VDD.n2262 0.3365
R5287 VDD.n2264 VDD.n2263 0.3365
R5288 VDD.n2265 VDD.n2264 0.3365
R5289 VDD.n2266 VDD.n2265 0.3365
R5290 VDD.n2267 VDD.n2266 0.3365
R5291 VDD.n2268 VDD.n2267 0.3365
R5292 VDD.n2269 VDD.n2268 0.3365
R5293 VDD.n2270 VDD.n2269 0.3365
R5294 VDD.n2314 VDD.n2313 0.3365
R5295 VDD.n1555 VDD.n1554 0.33575
R5296 VDD.n1657 VDD.n1656 0.33575
R5297 VDD.n1903 VDD.n1902 0.33575
R5298 VDD.n1405 VDD.n1404 0.335
R5299 VDD.n1358 VDD.n1357 0.33425
R5300 VDD.n1736 VDD.n1735 0.3335
R5301 VDD.n926 VDD.n925 0.33275
R5302 VDD.n2063 VDD.n2062 0.33275
R5303 VDD.n1401 VDD.n1400 0.3305
R5304 VDD.n1845 VDD.n1844 0.3305
R5305 VDD.n624 VDD.n623 0.3275
R5306 VDD.n1865 VDD.n1864 0.3275
R5307 VDD.n1972 VDD.n1971 0.3275
R5308 VDD.n284 VDD.n283 0.3275
R5309 VDD.n1677 VDD.n1676 0.32675
R5310 VDD.n1658 VDD.n1657 0.323
R5311 VDD.n1801 VDD.n1800 0.32225
R5312 VDD.n357 VDD.n356 0.32225
R5313 VDD.n2169 VDD.n2168 0.32225
R5314 VDD.n1458 VDD.n1457 0.3215
R5315 VDD.n1679 VDD.n1678 0.3215
R5316 VDD.n1869 VDD.n1868 0.3215
R5317 VDD.n1977 VDD.n1976 0.3215
R5318 VDD.n289 VDD.n288 0.3215
R5319 VDD.n1581 VDD.n1580 0.3185
R5320 VDD.n1864 VDD.n1863 0.3185
R5321 VDD.n1971 VDD.n1970 0.3185
R5322 VDD.n283 VDD.n282 0.3185
R5323 VDD.n1932 VDD.n1931 0.31475
R5324 VDD.n1562 VDD.n1561 0.314
R5325 VDD.n1549 VDD.n1548 0.314
R5326 VDD.n1536 VDD.n1535 0.314
R5327 VDD.n537 VDD.n536 0.314
R5328 VDD.n1363 VDD.n1362 0.314
R5329 VDD.n1841 VDD.n1840 0.314
R5330 VDD.n2041 VDD.n2040 0.314
R5331 VDD.n1567 VDD.n1566 0.3125
R5332 VDD.n1539 VDD.n1538 0.3125
R5333 VDD.n1617 VDD.n1616 0.3125
R5334 VDD.n452 VDD.n451 0.3125
R5335 VDD.n356 VDD.n355 0.3125
R5336 VDD.n1998 VDD.n1997 0.3125
R5337 VDD.n2010 VDD.n2009 0.3125
R5338 VDD.n2029 VDD.n2028 0.3125
R5339 VDD.n2061 VDD.n2060 0.3125
R5340 VDD.n2047 VDD.n2046 0.3125
R5341 VDD.n2316 VDD.n2315 0.3125
R5342 VDD.n1404 VDD.n1403 0.311
R5343 VDD.n1402 VDD.n1401 0.3095
R5344 VDD.n1291 VDD.n1290 0.30725
R5345 VDD.n1716 VDD.n1715 0.30725
R5346 VDD.n1505 VDD.n1504 0.3065
R5347 VDD.n1570 VDD.n1569 0.3065
R5348 VDD.n1537 VDD.n1536 0.3065
R5349 VDD.n1369 VDD.n1368 0.3065
R5350 VDD.n1593 VDD.n1592 0.3065
R5351 VDD.n1634 VDD.n1633 0.3065
R5352 VDD.n1300 VDD.n1299 0.3065
R5353 VDD.n1292 VDD.n1291 0.3065
R5354 VDD.n1725 VDD.n1724 0.3065
R5355 VDD.n1724 VDD.n1723 0.3065
R5356 VDD.n1698 VDD.n1697 0.3065
R5357 VDD.n1808 VDD.n1807 0.3065
R5358 VDD.n1102 VDD.n1101 0.3065
R5359 VDD.n1911 VDD.n1910 0.3065
R5360 VDD.n1909 VDD.n1908 0.3065
R5361 VDD.n1889 VDD.n1888 0.3065
R5362 VDD.n1931 VDD.n1930 0.3065
R5363 VDD.n1937 VDD.n1936 0.3065
R5364 VDD.n1945 VDD.n1944 0.3065
R5365 VDD.n2013 VDD.n2012 0.3065
R5366 VDD.n2057 VDD.n2056 0.3065
R5367 VDD.n2052 VDD.n2051 0.3065
R5368 VDD.n2049 VDD.n2048 0.3065
R5369 VDD.n2129 VDD.n2128 0.3065
R5370 VDD.n2167 VDD.n2166 0.3065
R5371 VDD.n2170 VDD.n2169 0.3065
R5372 VDD.n2319 VDD.n2318 0.3065
R5373 VDD.n144 VDD.n142 0.3055
R5374 VDD.n1410 VDD.n1409 0.30425
R5375 VDD.n1738 VDD.n1737 0.3035
R5376 VDD.n1734 VDD.n1733 0.3035
R5377 VDD.n1867 VDD.n1866 0.3035
R5378 VDD.n1974 VDD.n1973 0.3035
R5379 VDD.n286 VDD.n285 0.3035
R5380 VDD.n1360 VDD.n1359 0.3005
R5381 VDD.n174 VDD.n173 0.3005
R5382 VDD.n173 VDD.n172 0.3005
R5383 VDD.n172 VDD.n130 0.3005
R5384 VDD.n168 VDD.n130 0.3005
R5385 VDD.n168 VDD.n167 0.3005
R5386 VDD.n167 VDD.n166 0.3005
R5387 VDD.n163 VDD.n162 0.3005
R5388 VDD.n162 VDD.n161 0.3005
R5389 VDD.n161 VDD.n137 0.3005
R5390 VDD.n157 VDD.n137 0.3005
R5391 VDD.n157 VDD.n156 0.3005
R5392 VDD.n156 VDD.n155 0.3005
R5393 VDD.n152 VDD.n151 0.3005
R5394 VDD.n151 VDD.n150 0.3005
R5395 VDD.n150 VDD.n141 0.3005
R5396 VDD.n146 VDD.n141 0.3005
R5397 VDD.n146 VDD.n145 0.3005
R5398 VDD.n622 VDD.n621 0.298425
R5399 VDD.n1748 VDD.n1747 0.2975
R5400 VDD.n1856 VDD.n1855 0.29675
R5401 VDD.n1718 VDD.n1717 0.2945
R5402 VDD.n2012 VDD.n2011 0.2945
R5403 VDD.n1894 VDD.n1893 0.29375
R5404 VDD.n1668 VDD.n1667 0.29225
R5405 VDD.n1295 VDD.n1294 0.2915
R5406 VDD.n1467 VDD.n1466 0.2855
R5407 VDD.n1381 VDD.n1380 0.28475
R5408 VDD.n1563 VDD.n1562 0.284
R5409 VDD.n1313 VDD.n1312 0.2825
R5410 VDD.n1122 VDD.n1121 0.2825
R5411 VDD.n1984 VDD.n1983 0.2825
R5412 VDD.n942 VDD.n941 0.2825
R5413 VDD.n2160 VDD.n2159 0.2825
R5414 VDD.n2173 VDD.n2171 0.2825
R5415 VDD.n1307 VDD.n1306 0.28175
R5416 VDD.n1114 VDD.n1113 0.28175
R5417 VDD.n2171 VDD.n2170 0.28175
R5418 VDD.n120 VDD.n119 0.28175
R5419 VDD.n1483 VDD.n1481 0.281
R5420 VDD.n1429 VDD.n1428 0.2795
R5421 VDD.n1820 VDD.n1819 0.2795
R5422 VDD.n1891 VDD.n1890 0.2795
R5423 VDD.n1116 VDD.n1115 0.27875
R5424 VDD.n2131 VDD.n2130 0.278
R5425 VDD.n1729 VDD.n1728 0.2765
R5426 VDD.n1906 VDD.n1905 0.2765
R5427 VDD.n2138 VDD.n2137 0.2765
R5428 VDD.n2119 VDD.n2118 0.2765
R5429 VDD.n453 VDD.n452 0.27575
R5430 VDD.n1722 VDD.n1721 0.2735
R5431 VDD.n2008 VDD.n2007 0.2735
R5432 VDD.n2064 VDD.n2063 0.2735
R5433 VDD.n1656 VDD.n1655 0.272
R5434 VDD.n1626 VDD.n1625 0.27125
R5435 VDD.n454 VDD.n453 0.27125
R5436 VDD.n1638 VDD.n1637 0.2705
R5437 VDD.n1283 VDD.n1282 0.2705
R5438 VDD.n1455 VDD.n1454 0.2675
R5439 VDD.n1457 VDD.n1456 0.2675
R5440 VDD.n1720 VDD.n1719 0.2675
R5441 VDD.n1746 VDD.n1745 0.2675
R5442 VDD.n1773 VDD.n1772 0.2675
R5443 VDD.n1302 VDD.n1301 0.26675
R5444 VDD.n1895 VDD.n1894 0.266
R5445 VDD.n928 VDD.n927 0.266
R5446 VDD.n1644 VDD.n479 0.2645
R5447 VDD.n1571 VDD.n1570 0.263
R5448 VDD.n1500 VDD.n1499 0.26225
R5449 VDD.n7 VDD.n6 0.261581
R5450 VDD.n20 VDD.n19 0.261581
R5451 VDD.n32 VDD.n31 0.261581
R5452 VDD.n43 VDD.n42 0.261581
R5453 VDD.n55 VDD.n54 0.261581
R5454 VDD.n67 VDD.n66 0.261581
R5455 VDD.n79 VDD.n78 0.261581
R5456 VDD.n91 VDD.n90 0.261581
R5457 VDD.n1465 VDD.n1464 0.2615
R5458 VDD.n539 VDD.n538 0.2615
R5459 VDD.n448 VDD.n447 0.2615
R5460 VDD.n1797 VDD.n1796 0.2615
R5461 VDD.n353 VDD.n352 0.2615
R5462 VDD.n1943 VDD.n310 0.2615
R5463 VDD.n1899 VDD.n1898 0.26
R5464 VDD.n1751 VDD.n1750 0.25925
R5465 VDD.n2021 VDD.n2020 0.2585
R5466 VDD.n1633 VDD.n1632 0.25625
R5467 VDD.n1431 VDD.n1430 0.2555
R5468 VDD.n1662 VDD.n1661 0.2555
R5469 VDD.n1557 VDD.n1556 0.25475
R5470 VDD.n1526 VDD.n545 0.254
R5471 VDD.n1870 VDD.n1869 0.254
R5472 VDD.n2188 VDD.n2187 0.254
R5473 VDD.n144 VDD.n143 0.2535
R5474 VDD.n1481 VDD.n1480 0.25325
R5475 VDD.n626 VDD.n625 0.2525
R5476 VDD.n628 VDD.n627 0.2525
R5477 VDD.n630 VDD.n629 0.2525
R5478 VDD.n1446 VDD.n1445 0.2525
R5479 VDD.n1448 VDD.n1447 0.2525
R5480 VDD.n1450 VDD.n1449 0.2525
R5481 VDD.n1493 VDD.n1492 0.2525
R5482 VDD.n1377 VDD.n1376 0.2525
R5483 VDD.n1260 VDD.n1259 0.2525
R5484 VDD.n1258 VDD.n1257 0.2525
R5485 VDD.n1256 VDD.n1255 0.2525
R5486 VDD.n1254 VDD.n1253 0.2525
R5487 VDD.n1252 VDD.n1251 0.2525
R5488 VDD.n1250 VDD.n1249 0.2525
R5489 VDD.n1327 VDD.n1326 0.2525
R5490 VDD.n1325 VDD.n1324 0.2525
R5491 VDD.n1323 VDD.n1322 0.2525
R5492 VDD.n1321 VDD.n1320 0.2525
R5493 VDD.n1319 VDD.n1318 0.2525
R5494 VDD.n1317 VDD.n1316 0.2525
R5495 VDD.n1315 VDD.n1314 0.2525
R5496 VDD.n1311 VDD.n1310 0.2525
R5497 VDD.n1219 VDD.n1218 0.2525
R5498 VDD.n1217 VDD.n1216 0.2525
R5499 VDD.n1215 VDD.n1214 0.2525
R5500 VDD.n1213 VDD.n1212 0.2525
R5501 VDD.n1211 VDD.n1210 0.2525
R5502 VDD.n1209 VDD.n1208 0.2525
R5503 VDD.n1242 VDD.n1241 0.2525
R5504 VDD.n1240 VDD.n1239 0.2525
R5505 VDD.n1238 VDD.n1237 0.2525
R5506 VDD.n1236 VDD.n1235 0.2525
R5507 VDD.n1234 VDD.n1233 0.2525
R5508 VDD.n1232 VDD.n1231 0.2525
R5509 VDD.n1230 VDD.n1229 0.2525
R5510 VDD.n1228 VDD.n1227 0.2525
R5511 VDD.n1173 VDD.n1172 0.2525
R5512 VDD.n1171 VDD.n1170 0.2525
R5513 VDD.n1169 VDD.n1168 0.2525
R5514 VDD.n1167 VDD.n1166 0.2525
R5515 VDD.n1165 VDD.n1164 0.2525
R5516 VDD.n1163 VDD.n1162 0.2525
R5517 VDD.n1822 VDD.n1821 0.2525
R5518 VDD.n1818 VDD.n1817 0.2525
R5519 VDD.n1816 VDD.n1815 0.2525
R5520 VDD.n1814 VDD.n1813 0.2525
R5521 VDD.n1812 VDD.n1811 0.2525
R5522 VDD.n1087 VDD.n1086 0.2525
R5523 VDD.n1085 VDD.n1084 0.2525
R5524 VDD.n1083 VDD.n1082 0.2525
R5525 VDD.n1081 VDD.n1080 0.2525
R5526 VDD.n1079 VDD.n1078 0.2525
R5527 VDD.n1077 VDD.n1076 0.2525
R5528 VDD.n1155 VDD.n1154 0.2525
R5529 VDD.n1153 VDD.n1152 0.2525
R5530 VDD.n1151 VDD.n1150 0.2525
R5531 VDD.n1149 VDD.n1148 0.2525
R5532 VDD.n1147 VDD.n1146 0.2525
R5533 VDD.n1145 VDD.n1144 0.2525
R5534 VDD.n1143 VDD.n1142 0.2525
R5535 VDD.n1141 VDD.n1140 0.2525
R5536 VDD.n1137 VDD.n1136 0.2525
R5537 VDD.n1135 VDD.n1134 0.2525
R5538 VDD.n1133 VDD.n1132 0.2525
R5539 VDD.n1131 VDD.n1130 0.2525
R5540 VDD.n1129 VDD.n1128 0.2525
R5541 VDD.n1124 VDD.n1123 0.2525
R5542 VDD.n1040 VDD.n1039 0.2525
R5543 VDD.n1038 VDD.n1037 0.2525
R5544 VDD.n1036 VDD.n1035 0.2525
R5545 VDD.n1034 VDD.n1033 0.2525
R5546 VDD.n1032 VDD.n1031 0.2525
R5547 VDD.n1030 VDD.n1029 0.2525
R5548 VDD.n1069 VDD.n1068 0.2525
R5549 VDD.n1067 VDD.n1066 0.2525
R5550 VDD.n1065 VDD.n1064 0.2525
R5551 VDD.n1063 VDD.n1062 0.2525
R5552 VDD.n1061 VDD.n1060 0.2525
R5553 VDD.n1059 VDD.n1058 0.2525
R5554 VDD.n1057 VDD.n1056 0.2525
R5555 VDD.n1055 VDD.n1054 0.2525
R5556 VDD.n1051 VDD.n1050 0.2525
R5557 VDD.n1049 VDD.n1048 0.2525
R5558 VDD.n1047 VDD.n1046 0.2525
R5559 VDD.n1045 VDD.n1044 0.2525
R5560 VDD.n1043 VDD.n1042 0.2525
R5561 VDD.n1917 VDD.n1916 0.2525
R5562 VDD.n1915 VDD.n1914 0.2525
R5563 VDD.n993 VDD.n992 0.2525
R5564 VDD.n991 VDD.n990 0.2525
R5565 VDD.n989 VDD.n988 0.2525
R5566 VDD.n987 VDD.n986 0.2525
R5567 VDD.n985 VDD.n984 0.2525
R5568 VDD.n983 VDD.n982 0.2525
R5569 VDD.n1022 VDD.n1021 0.2525
R5570 VDD.n1020 VDD.n1019 0.2525
R5571 VDD.n1018 VDD.n1017 0.2525
R5572 VDD.n1016 VDD.n1015 0.2525
R5573 VDD.n1014 VDD.n1013 0.2525
R5574 VDD.n1012 VDD.n1011 0.2525
R5575 VDD.n1010 VDD.n1009 0.2525
R5576 VDD.n1008 VDD.n1007 0.2525
R5577 VDD.n1004 VDD.n1003 0.2525
R5578 VDD.n1002 VDD.n1001 0.2525
R5579 VDD.n1000 VDD.n999 0.2525
R5580 VDD.n998 VDD.n997 0.2525
R5581 VDD.n996 VDD.n995 0.2525
R5582 VDD.n1925 VDD.n1924 0.2525
R5583 VDD.n1927 VDD.n1926 0.2525
R5584 VDD.n913 VDD.n912 0.2525
R5585 VDD.n911 VDD.n910 0.2525
R5586 VDD.n909 VDD.n908 0.2525
R5587 VDD.n907 VDD.n906 0.2525
R5588 VDD.n905 VDD.n904 0.2525
R5589 VDD.n903 VDD.n902 0.2525
R5590 VDD.n975 VDD.n974 0.2525
R5591 VDD.n973 VDD.n972 0.2525
R5592 VDD.n971 VDD.n970 0.2525
R5593 VDD.n969 VDD.n968 0.2525
R5594 VDD.n967 VDD.n966 0.2525
R5595 VDD.n965 VDD.n964 0.2525
R5596 VDD.n963 VDD.n962 0.2525
R5597 VDD.n961 VDD.n960 0.2525
R5598 VDD.n957 VDD.n956 0.2525
R5599 VDD.n955 VDD.n954 0.2525
R5600 VDD.n953 VDD.n952 0.2525
R5601 VDD.n951 VDD.n950 0.2525
R5602 VDD.n949 VDD.n948 0.2525
R5603 VDD.n944 VDD.n943 0.2525
R5604 VDD.n939 VDD.n938 0.2525
R5605 VDD.n937 VDD.n936 0.2525
R5606 VDD.n935 VDD.n934 0.2525
R5607 VDD.n933 VDD.n932 0.2525
R5608 VDD.n866 VDD.n865 0.2525
R5609 VDD.n864 VDD.n863 0.2525
R5610 VDD.n862 VDD.n861 0.2525
R5611 VDD.n860 VDD.n859 0.2525
R5612 VDD.n858 VDD.n857 0.2525
R5613 VDD.n856 VDD.n855 0.2525
R5614 VDD.n895 VDD.n894 0.2525
R5615 VDD.n893 VDD.n892 0.2525
R5616 VDD.n891 VDD.n890 0.2525
R5617 VDD.n889 VDD.n888 0.2525
R5618 VDD.n887 VDD.n886 0.2525
R5619 VDD.n885 VDD.n884 0.2525
R5620 VDD.n883 VDD.n882 0.2525
R5621 VDD.n881 VDD.n880 0.2525
R5622 VDD.n877 VDD.n876 0.2525
R5623 VDD.n875 VDD.n874 0.2525
R5624 VDD.n873 VDD.n872 0.2525
R5625 VDD.n871 VDD.n870 0.2525
R5626 VDD.n869 VDD.n868 0.2525
R5627 VDD.n2078 VDD.n2077 0.2525
R5628 VDD.n2076 VDD.n2075 0.2525
R5629 VDD.n819 VDD.n818 0.2525
R5630 VDD.n817 VDD.n816 0.2525
R5631 VDD.n815 VDD.n814 0.2525
R5632 VDD.n813 VDD.n812 0.2525
R5633 VDD.n811 VDD.n810 0.2525
R5634 VDD.n809 VDD.n808 0.2525
R5635 VDD.n848 VDD.n847 0.2525
R5636 VDD.n846 VDD.n845 0.2525
R5637 VDD.n844 VDD.n843 0.2525
R5638 VDD.n842 VDD.n841 0.2525
R5639 VDD.n840 VDD.n839 0.2525
R5640 VDD.n838 VDD.n837 0.2525
R5641 VDD.n836 VDD.n835 0.2525
R5642 VDD.n834 VDD.n833 0.2525
R5643 VDD.n830 VDD.n829 0.2525
R5644 VDD.n828 VDD.n827 0.2525
R5645 VDD.n826 VDD.n825 0.2525
R5646 VDD.n824 VDD.n823 0.2525
R5647 VDD.n822 VDD.n821 0.2525
R5648 VDD.n2086 VDD.n2085 0.2525
R5649 VDD.n2088 VDD.n2087 0.2525
R5650 VDD.n740 VDD.n739 0.2525
R5651 VDD.n738 VDD.n737 0.2525
R5652 VDD.n736 VDD.n735 0.2525
R5653 VDD.n734 VDD.n733 0.2525
R5654 VDD.n732 VDD.n731 0.2525
R5655 VDD.n730 VDD.n729 0.2525
R5656 VDD.n801 VDD.n800 0.2525
R5657 VDD.n799 VDD.n798 0.2525
R5658 VDD.n797 VDD.n796 0.2525
R5659 VDD.n795 VDD.n794 0.2525
R5660 VDD.n793 VDD.n792 0.2525
R5661 VDD.n791 VDD.n790 0.2525
R5662 VDD.n789 VDD.n788 0.2525
R5663 VDD.n787 VDD.n786 0.2525
R5664 VDD.n783 VDD.n782 0.2525
R5665 VDD.n781 VDD.n780 0.2525
R5666 VDD.n779 VDD.n778 0.2525
R5667 VDD.n777 VDD.n776 0.2525
R5668 VDD.n775 VDD.n774 0.2525
R5669 VDD.n770 VDD.n769 0.2525
R5670 VDD.n768 VDD.n767 0.2525
R5671 VDD.n764 VDD.n763 0.2525
R5672 VDD.n762 VDD.n761 0.2525
R5673 VDD.n760 VDD.n759 0.2525
R5674 VDD.n758 VDD.n757 0.2525
R5675 VDD.n756 VDD.n755 0.2525
R5676 VDD.n754 VDD.n753 0.2525
R5677 VDD.n752 VDD.n751 0.2525
R5678 VDD.n750 VDD.n749 0.2525
R5679 VDD.n746 VDD.n745 0.2525
R5680 VDD.n744 VDD.n743 0.2525
R5681 VDD.n742 VDD.n239 0.2525
R5682 VDD.n2154 VDD.n2153 0.2525
R5683 VDD.n2156 VDD.n2155 0.2525
R5684 VDD.n2162 VDD.n2161 0.2525
R5685 VDD.n2165 VDD.n2164 0.2525
R5686 VDD.n693 VDD.n692 0.2525
R5687 VDD.n691 VDD.n690 0.2525
R5688 VDD.n689 VDD.n688 0.2525
R5689 VDD.n687 VDD.n686 0.2525
R5690 VDD.n685 VDD.n684 0.2525
R5691 VDD.n683 VDD.n682 0.2525
R5692 VDD.n722 VDD.n721 0.2525
R5693 VDD.n720 VDD.n719 0.2525
R5694 VDD.n718 VDD.n717 0.2525
R5695 VDD.n716 VDD.n715 0.2525
R5696 VDD.n714 VDD.n713 0.2525
R5697 VDD.n712 VDD.n711 0.2525
R5698 VDD.n710 VDD.n709 0.2525
R5699 VDD.n708 VDD.n707 0.2525
R5700 VDD.n704 VDD.n703 0.2525
R5701 VDD.n702 VDD.n701 0.2525
R5702 VDD.n700 VDD.n699 0.2525
R5703 VDD.n698 VDD.n697 0.2525
R5704 VDD.n696 VDD.n695 0.2525
R5705 VDD.n2250 VDD.n2249 0.2525
R5706 VDD.n2248 VDD.n2247 0.2525
R5707 VDD.n2244 VDD.n2243 0.2525
R5708 VDD.n2242 VDD.n2241 0.2525
R5709 VDD.n2240 VDD.n2239 0.2525
R5710 VDD.n2238 VDD.n2237 0.2525
R5711 VDD.n2236 VDD.n2235 0.2525
R5712 VDD.n2234 VDD.n2233 0.2525
R5713 VDD.n2232 VDD.n2231 0.2525
R5714 VDD.n2230 VDD.n2229 0.2525
R5715 VDD.n2226 VDD.n2225 0.2525
R5716 VDD.n2224 VDD.n2223 0.2525
R5717 VDD.n2222 VDD.n2221 0.2525
R5718 VDD.n2217 VDD.n2216 0.2525
R5719 VDD.n2215 VDD.n2214 0.2525
R5720 VDD.n2213 VDD.n2212 0.2525
R5721 VDD.n2211 VDD.n2210 0.2525
R5722 VDD.n2199 VDD.n2198 0.2525
R5723 VDD.n2197 VDD.n2196 0.2525
R5724 VDD.n2195 VDD.n2194 0.2525
R5725 VDD.n2317 VDD.n2316 0.2525
R5726 VDD.n1309 VDD.n1308 0.25175
R5727 VDD.n1999 VDD.n1998 0.251
R5728 VDD.n2192 VDD.n2191 0.251
R5729 VDD.n1673 VDD.n1672 0.2495
R5730 VDD.n1690 VDD.n1689 0.24875
R5731 VDD.n1934 VDD.n1933 0.24875
R5732 VDD.n200 VDD.n199 0.248188
R5733 VDD.n1280 VDD.n1279 0.248
R5734 VDD.n2124 VDD.n2123 0.248
R5735 VDD.n1991 VDD.n1990 0.24725
R5736 VDD.n1276 VDD.n1275 0.2465
R5737 VDD.n1554 VDD.n1553 0.24425
R5738 VDD.n1511 VDD.n1510 0.2435
R5739 VDD.n1862 VDD.n1861 0.2435
R5740 VDD.n1969 VDD.n1968 0.2435
R5741 VDD.n281 VDD.n280 0.2435
R5742 VDD.n1640 VDD.n1639 0.242
R5743 VDD.n1654 VDD.n1653 0.2405
R5744 VDD.n1809 VDD.n1808 0.2405
R5745 VDD.n1588 VDD.n1587 0.23975
R5746 VDD.n2149 VDD.n243 0.239
R5747 VDD.n455 VDD.n454 0.23825
R5748 VDD.n1938 VDD.n1937 0.23825
R5749 VDD.n632 VDD.n631 0.2375
R5750 VDD.n1444 VDD.n1443 0.2375
R5751 VDD.n1543 VDD.n1542 0.2375
R5752 VDD.n1831 VDD.n1830 0.2375
R5753 VDD.n1596 VDD.n1589 0.23675
R5754 VDD.n2336 VDD.n109 0.235598
R5755 VDD.n1800 VDD.n1799 0.2345
R5756 VDD.n1112 VDD.n1111 0.2345
R5757 VDD.n2219 VDD.n2218 0.233
R5758 VDD.n1417 VDD.n1373 0.23
R5759 VDD.n1371 VDD.n1333 0.23
R5760 VDD.n1331 VDD.n1248 0.23
R5761 VDD.n1246 VDD.n1207 0.23
R5762 VDD.n1205 VDD.n1161 0.23
R5763 VDD.n1159 VDD.n1075 0.23
R5764 VDD.n1073 VDD.n1028 0.23
R5765 VDD.n1026 VDD.n981 0.23
R5766 VDD.n979 VDD.n901 0.23
R5767 VDD.n899 VDD.n854 0.23
R5768 VDD.n2039 VDD.n2038 0.23
R5769 VDD.n852 VDD.n807 0.23
R5770 VDD.n2140 VDD.n2139 0.23
R5771 VDD.n805 VDD.n728 0.23
R5772 VDD.n726 VDD.n681 0.23
R5773 VDD.n1434 VDD.n1433 0.2285
R5774 VDD.n1367 VDD.n1366 0.2285
R5775 VDD.n1730 VDD.n1729 0.2285
R5776 VDD.n1699 VDD.n1698 0.2285
R5777 VDD.n1907 VDD.n1906 0.2285
R5778 VDD.n1840 VDD.n1839 0.22775
R5779 VDD.n2003 VDD.n2002 0.22775
R5780 VDD.n2143 VDD.n2142 0.22775
R5781 VDD.n1627 VDD.n1626 0.22625
R5782 VDD.n1288 VDD.n1287 0.22625
R5783 VDD.n1892 VDD.n1891 0.2255
R5784 VDD.n1299 VDD.n1298 0.22325
R5785 VDD.n1329 VDD.n1328 0.2225
R5786 VDD.n1226 VDD.n1225 0.2225
R5787 VDD.n1203 VDD.n1202 0.2225
R5788 VDD.n1139 VDD.n1138 0.2225
R5789 VDD.n1913 VDD.n1912 0.2225
R5790 VDD.n1878 VDD.n1877 0.2225
R5791 VDD.n1929 VDD.n1928 0.2225
R5792 VDD.n1993 VDD.n1992 0.2225
R5793 VDD.n959 VDD.n958 0.2225
R5794 VDD.n2006 VDD.n2005 0.2225
R5795 VDD.n2074 VDD.n2073 0.2225
R5796 VDD.n2090 VDD.n2089 0.2225
R5797 VDD.n748 VDD.n747 0.2225
R5798 VDD.n2209 VDD.n2208 0.2225
R5799 VDD.n2193 VDD.n2192 0.2225
R5800 VDD.n1304 VDD.n1303 0.221
R5801 VDD.n1462 VDD.n1461 0.2195
R5802 VDD.n1285 VDD.n1284 0.2195
R5803 VDD.n1933 VDD.n1932 0.2195
R5804 VDD.n1624 VDD.n1623 0.21875
R5805 VDD.n1807 VDD.n1806 0.21875
R5806 VDD.n1877 VDD.n1876 0.21875
R5807 VDD.n1983 VDD.n1982 0.21875
R5808 VDD.n2058 VDD.n2057 0.21875
R5809 VDD.n2038 VDD.n2037 0.21875
R5810 VDD.n1763 VDD.n1762 0.2165
R5811 VDD.n1765 VDD.n1764 0.2165
R5812 VDD.n1948 VDD.n1947 0.2165
R5813 VDD.n541 VDD.n540 0.215
R5814 VDD.n1648 VDD.n1647 0.21425
R5815 VDD.n163 VDD.n135 0.21425
R5816 VDD.n1440 VDD.n1439 0.2135
R5817 VDD.n1646 VDD.n1645 0.2135
R5818 VDD.n1705 VDD.n1704 0.2135
R5819 VDD.n1703 VDD.n1702 0.2135
R5820 VDD.n1701 VDD.n1700 0.2135
R5821 VDD.n1689 VDD.n1688 0.2135
R5822 VDD.n1833 VDD.n1832 0.2135
R5823 VDD.n1740 VDD.n1739 0.212
R5824 VDD.n1744 VDD.n1743 0.212
R5825 VDD.n1126 VDD.n1125 0.212
R5826 VDD.n946 VDD.n945 0.212
R5827 VDD.n2256 VDD.n2255 0.212
R5828 VDD VDD.n0 0.211771
R5829 VDD.n1829 VDD.n1828 0.21125
R5830 VDD.t1425 VDD.t415 0.210232
R5831 VDD.n1362 VDD.n1361 0.20975
R5832 VDD.n1534 VDD.n1533 0.209
R5833 VDD.n1710 VDD.n1709 0.209
R5834 VDD.n1497 VDD.n1496 0.20825
R5835 VDD.n544 VDD.n543 0.20825
R5836 VDD.n1474 VDD.n1473 0.2075
R5837 VDD.n1774 VDD.n1773 0.2075
R5838 VDD.n1109 VDD.n1108 0.2075
R5839 VDD.n1660 VDD.n1659 0.206
R5840 VDD.n1178 VDD.n405 0.20525
R5841 VDD.n1282 VDD.n1281 0.2045
R5842 VDD.n1713 VDD.n1712 0.20225
R5843 VDD.n2121 VDD.n2120 0.2015
R5844 VDD.n1635 VDD.n1634 0.20075
R5845 VDD.n1650 VDD.n1649 0.19925
R5846 VDD.n1407 VDD.n1406 0.1985
R5847 VDD.n1187 VDD.n1186 0.1985
R5848 VDD.n659 VDD.n658 0.1985
R5849 VDD.n2261 VDD.n2260 0.1985
R5850 VDD.n2322 VDD.n2321 0.1985
R5851 VDD.n2305 VDD.n2304 0.1985
R5852 VDD.n1631 VDD.n1630 0.19625
R5853 VDD.n2048 VDD.n2047 0.19625
R5854 VDD.n1485 VDD.n1484 0.1955
R5855 VDD.n1504 VDD.n1503 0.19475
R5856 VDD.n1384 VDD.n1383 0.19475
R5857 VDD.n1281 VDD.n1280 0.194
R5858 VDD.n1491 VDD.n1490 0.1925
R5859 VDD.n1879 VDD.n1878 0.191
R5860 VDD.n2132 VDD.n2131 0.191
R5861 VDD.n1755 VDD.n1754 0.1895
R5862 VDD.n1757 VDD.n1756 0.1895
R5863 VDD.n1759 VDD.n1758 0.1895
R5864 VDD.n1761 VDD.n1760 0.1895
R5865 VDD.n1522 VDD.n1521 0.1835
R5866 VDD.n536 VDD.n535 0.1835
R5867 VDD.n2040 VDD.n2039 0.1835
R5868 VDD.n2185 VDD.n2184 0.1835
R5869 VDD.n2183 VDD.n2182 0.1835
R5870 VDD.n2181 VDD.n2180 0.1835
R5871 VDD.n2179 VDD.n2178 0.1835
R5872 VDD.n2177 VDD.n2176 0.1835
R5873 VDD.n2297 VDD.n2296 0.1835
R5874 VDD.n2295 VDD.n2294 0.1835
R5875 VDD.n2293 VDD.n2292 0.1835
R5876 VDD.n2291 VDD.n2290 0.1835
R5877 VDD.n2289 VDD.n2288 0.1835
R5878 VDD.n1902 VDD.n1901 0.18275
R5879 VDD.n1421 VDD.n1420 0.182
R5880 VDD.n1827 VDD.n1826 0.18125
R5881 VDD.n1839 VDD.n1838 0.18125
R5882 VDD.n1671 VDD.n1670 0.1775
R5883 VDD.n1771 VDD.n1770 0.1775
R5884 VDD.n155 VDD.n139 0.17675
R5885 VDD.n1479 VDD.n1478 0.17525
R5886 VDD.n1413 VDD.n1412 0.1745
R5887 VDD.n1629 VDD.n1628 0.1745
R5888 VDD.n1422 VDD.n1421 0.17375
R5889 VDD.n1470 VDD.n1469 0.17375
R5890 VDD.n1487 VDD.n1486 0.1715
R5891 VDD.n1107 VDD.n1106 0.1715
R5892 VDD.n1427 VDD.n1426 0.16925
R5893 VDD.n1437 VDD.n1436 0.1685
R5894 VDD.n1520 VDD.n1519 0.1685
R5895 VDD.n1519 VDD.n1518 0.1685
R5896 VDD.n1518 VDD.n1517 0.1685
R5897 VDD.n1517 VDD.n1516 0.1685
R5898 VDD.n1516 VDD.n1515 0.1685
R5899 VDD.n1515 VDD.n1514 0.1685
R5900 VDD.n1514 VDD.n1513 0.1685
R5901 VDD.n1513 VDD.n1512 0.1685
R5902 VDD.n1512 VDD.n1511 0.1685
R5903 VDD.n1408 VDD.n1407 0.1685
R5904 VDD.n1613 VDD.n1612 0.1685
R5905 VDD.n1202 VDD.n1201 0.1685
R5906 VDD.n1201 VDD.n1200 0.1685
R5907 VDD.n1200 VDD.n1199 0.1685
R5908 VDD.n1199 VDD.n1198 0.1685
R5909 VDD.n1198 VDD.n1197 0.1685
R5910 VDD.n1197 VDD.n1196 0.1685
R5911 VDD.n1196 VDD.n1195 0.1685
R5912 VDD.n1195 VDD.n1194 0.1685
R5913 VDD.n1194 VDD.n1193 0.1685
R5914 VDD.n1193 VDD.n1192 0.1685
R5915 VDD.n1192 VDD.n1191 0.1685
R5916 VDD.n1191 VDD.n1190 0.1685
R5917 VDD.n1190 VDD.n1189 0.1685
R5918 VDD.n1189 VDD.n1188 0.1685
R5919 VDD.n1188 VDD.n1187 0.1685
R5920 VDD.n1185 VDD.n1184 0.1685
R5921 VDD.n1184 VDD.n1183 0.1685
R5922 VDD.n1183 VDD.n1182 0.1685
R5923 VDD.n2067 VDD.n2066 0.1685
R5924 VDD.n2066 VDD.n2065 0.1685
R5925 VDD.n2187 VDD.n2186 0.1685
R5926 VDD.n2208 VDD.n2207 0.1685
R5927 VDD.n2207 VDD.n2206 0.1685
R5928 VDD.n2206 VDD.n2205 0.1685
R5929 VDD.n2205 VDD.n2204 0.1685
R5930 VDD.n2204 VDD.n2203 0.1685
R5931 VDD.n2203 VDD.n2202 0.1685
R5932 VDD.n2202 VDD.n2201 0.1685
R5933 VDD.n2201 VDD.n2200 0.1685
R5934 VDD.n649 VDD.n648 0.1685
R5935 VDD.n648 VDD.n647 0.1685
R5936 VDD.n647 VDD.n646 0.1685
R5937 VDD.n646 VDD.n645 0.1685
R5938 VDD.n645 VDD.n644 0.1685
R5939 VDD.n644 VDD.n643 0.1685
R5940 VDD.n643 VDD.n642 0.1685
R5941 VDD.n642 VDD.n641 0.1685
R5942 VDD.n641 VDD.n640 0.1685
R5943 VDD.n640 VDD.n639 0.1685
R5944 VDD.n639 VDD.n638 0.1685
R5945 VDD.n638 VDD.n637 0.1685
R5946 VDD.n674 VDD.n673 0.1685
R5947 VDD.n673 VDD.n672 0.1685
R5948 VDD.n672 VDD.n671 0.1685
R5949 VDD.n671 VDD.n670 0.1685
R5950 VDD.n670 VDD.n669 0.1685
R5951 VDD.n669 VDD.n668 0.1685
R5952 VDD.n668 VDD.n667 0.1685
R5953 VDD.n667 VDD.n666 0.1685
R5954 VDD.n666 VDD.n665 0.1685
R5955 VDD.n665 VDD.n664 0.1685
R5956 VDD.n664 VDD.n663 0.1685
R5957 VDD.n663 VDD.n662 0.1685
R5958 VDD.n662 VDD.n661 0.1685
R5959 VDD.n661 VDD.n660 0.1685
R5960 VDD.n660 VDD.n659 0.1685
R5961 VDD.n2275 VDD.n2274 0.1685
R5962 VDD.n2274 VDD.n2273 0.1685
R5963 VDD.n2273 VDD.n2272 0.1685
R5964 VDD.n2272 VDD.n2271 0.1685
R5965 VDD.n2271 VDD.n217 0.1685
R5966 VDD.n2330 VDD.n2329 0.1685
R5967 VDD.n2329 VDD.n2328 0.1685
R5968 VDD.n2328 VDD.n2327 0.1685
R5969 VDD.n2327 VDD.n2326 0.1685
R5970 VDD.n2326 VDD.n2325 0.1685
R5971 VDD.n2325 VDD.n2324 0.1685
R5972 VDD.n2324 VDD.n2323 0.1685
R5973 VDD.n2323 VDD.n2322 0.1685
R5974 VDD.n2313 VDD.n2312 0.1685
R5975 VDD.n2312 VDD.n2311 0.1685
R5976 VDD.n2311 VDD.n2310 0.1685
R5977 VDD.n2310 VDD.n2309 0.1685
R5978 VDD.n2309 VDD.n2308 0.1685
R5979 VDD.n2308 VDD.n2307 0.1685
R5980 VDD.n2307 VDD.n2306 0.1685
R5981 VDD.n2306 VDD.n2305 0.1685
R5982 VDD.n2303 VDD.n2302 0.1685
R5983 VDD.n2300 VDD.n2299 0.1685
R5984 VDD.n2299 VDD.n2298 0.1685
R5985 VDD.n1641 VDD.n1640 0.167
R5986 VDD.n1488 VDD.n1487 0.1655
R5987 VDD.n2044 VDD.n2043 0.164
R5988 VDD.n1469 VDD.n1468 0.16325
R5989 VDD.n1592 VDD.n1591 0.16325
R5990 VDD.n1552 VDD.n1551 0.16175
R5991 VDD.n1620 VDD.n1619 0.16025
R5992 VDD.n1685 VDD.n455 0.16025
R5993 VDD.n1803 VDD.n1802 0.16025
R5994 VDD.n1873 VDD.n358 0.16025
R5995 VDD.n1979 VDD.n1978 0.16025
R5996 VDD.n2034 VDD.n290 0.16025
R5997 VDD.n1672 VDD.n1671 0.1595
R5998 VDD.n1708 VDD.n1707 0.1595
R5999 VDD.n1706 VDD.n1705 0.1595
R6000 VDD.n1770 VDD.n381 0.1595
R6001 VDD.n2050 VDD.n2049 0.15875
R6002 VDD.n2059 VDD.n2058 0.15575
R6003 VDD.n1530 VDD.n1529 0.15425
R6004 VDD.n1436 VDD.n1435 0.1535
R6005 VDD.n1521 VDD.n1520 0.1535
R6006 VDD.n535 VDD.n534 0.1535
R6007 VDD.n1796 VDD.n1795 0.1535
R6008 VDD.n2186 VDD.n2185 0.1535
R6009 VDD.n2184 VDD.n2183 0.1535
R6010 VDD.n2182 VDD.n2181 0.1535
R6011 VDD.n2180 VDD.n2179 0.1535
R6012 VDD.n2178 VDD.n2177 0.1535
R6013 VDD.n2176 VDD.n2175 0.1535
R6014 VDD.n2298 VDD.n2297 0.1535
R6015 VDD.n2296 VDD.n2295 0.1535
R6016 VDD.n2294 VDD.n2293 0.1535
R6017 VDD.n2292 VDD.n2291 0.1535
R6018 VDD.n2290 VDD.n2289 0.1535
R6019 VDD.n2288 VDD.n2287 0.1535
R6020 VDD.n1556 VDD.n1555 0.1505
R6021 VDD.n1293 VDD.n1292 0.1505
R6022 VDD.n1531 VDD.n1530 0.149
R6023 VDD.n2331 VDD.n2330 0.149
R6024 VDD.n1461 VDD.n1460 0.1475
R6025 VDD.n1707 VDD.n1706 0.1475
R6026 VDD.n1754 VDD.n1753 0.1475
R6027 VDD.n1756 VDD.n1755 0.1475
R6028 VDD.n1758 VDD.n1757 0.1475
R6029 VDD.n1760 VDD.n1759 0.1475
R6030 VDD.n1762 VDD.n1761 0.1475
R6031 VDD.n1686 VDD.n1685 0.14675
R6032 VDD.n1980 VDD.n1979 0.14675
R6033 VDD.n1420 VDD.n634 0.146
R6034 VDD.n1545 VDD.n1544 0.146
R6035 VDD.n1625 VDD.n1624 0.146
R6036 VDD.n1565 VDD.n1564 0.14525
R6037 VDD.n1944 VDD.n1943 0.14525
R6038 VDD.n1490 VDD.n1489 0.1445
R6039 VDD.n1621 VDD.n1620 0.1445
R6040 VDD.n1995 VDD.n1994 0.1445
R6041 VDD.n1442 VDD.n1441 0.14375
R6042 VDD.n1569 VDD.n1568 0.14375
R6043 VDD.n1651 VDD.n1650 0.14375
R6044 VDD.n2141 VDD.n2140 0.14375
R6045 VDD.n117 VDD.n116 0.143273
R6046 VDD.n1383 VDD.n1382 0.14225
R6047 VDD.n1753 VDD.n1752 0.14225
R6048 VDD.n1486 VDD.n1485 0.1415
R6049 VDD.n1719 VDD.n1718 0.1415
R6050 VDD.n186 VDD.n185 0.141125
R6051 VDD.n1804 VDD.n1803 0.14075
R6052 VDD.n1874 VDD.n1873 0.14075
R6053 VDD.n1523 VDD.n548 0.14
R6054 VDD.n1616 VDD.n1615 0.14
R6055 VDD.n179 VDD.n178 0.139447
R6056 VDD.n650 VDD.n649 0.139327
R6057 VDD.n1425 VDD.n1424 0.1385
R6058 VDD.n1476 VDD.n1475 0.1385
R6059 VDD.n1494 VDD.n1493 0.1385
R6060 VDD.n1507 VDD.n1506 0.1385
R6061 VDD.n1596 VDD.n1595 0.1385
R6062 VDD.n1244 VDD.n1243 0.1385
R6063 VDD.n1186 VDD.n1185 0.1385
R6064 VDD.n1824 VDD.n1823 0.1385
R6065 VDD.n1157 VDD.n1156 0.1385
R6066 VDD.n1071 VDD.n1070 0.1385
R6067 VDD.n1053 VDD.n1052 0.1385
R6068 VDD.n1024 VDD.n1023 0.1385
R6069 VDD.n1006 VDD.n1005 0.1385
R6070 VDD.n977 VDD.n976 0.1385
R6071 VDD.n897 VDD.n896 0.1385
R6072 VDD.n879 VDD.n878 0.1385
R6073 VDD.n850 VDD.n849 0.1385
R6074 VDD.n832 VDD.n831 0.1385
R6075 VDD.n803 VDD.n802 0.1385
R6076 VDD.n785 VDD.n784 0.1385
R6077 VDD.n766 VDD.n765 0.1385
R6078 VDD.n724 VDD.n723 0.1385
R6079 VDD.n706 VDD.n705 0.1385
R6080 VDD.n2246 VDD.n2245 0.1385
R6081 VDD.n2228 VDD.n2227 0.1385
R6082 VDD.n678 VDD.n677 0.1385
R6083 VDD.n675 VDD.n674 0.1385
R6084 VDD.n658 VDD.n657 0.1385
R6085 VDD.n2260 VDD.n2259 0.1385
R6086 VDD.n2262 VDD.n2261 0.1385
R6087 VDD.n2276 VDD.n2275 0.1385
R6088 VDD.n2321 VDD.n2320 0.1385
R6089 VDD.n2304 VDD.n2303 0.1385
R6090 VDD.n1417 VDD.n1416 0.137
R6091 VDD.n2026 VDD.n2025 0.137
R6092 VDD.n679 VDD.n678 0.137
R6093 VDD.n1352 VDD.n498 0.13625
R6094 VDD.n1731 VDD.n1730 0.1355
R6095 VDD.n449 VDD.n448 0.1355
R6096 VDD.n1452 VDD.n1451 0.134
R6097 VDD.n1870 VDD.n361 0.134
R6098 VDD.n1471 VDD.n1470 0.13325
R6099 VDD.n1682 VDD.n458 0.13325
R6100 VDD.n8 VDD.n7 0.131992
R6101 VDD.n21 VDD.n20 0.131992
R6102 VDD.n33 VDD.n32 0.131992
R6103 VDD.n44 VDD.n43 0.131992
R6104 VDD.n56 VDD.n55 0.131992
R6105 VDD.n68 VDD.n67 0.131992
R6106 VDD.n80 VDD.n79 0.131992
R6107 VDD.n92 VDD.n91 0.131992
R6108 VDD.n1480 VDD.n1479 0.13175
R6109 VDD.n1548 VDD.n1547 0.13175
R6110 VDD.n113 VDD.n112 0.131409
R6111 VDD.n118 VDD.n117 0.131409
R6112 VDD.n1443 VDD.n1442 0.1295
R6113 VDD.n1810 VDD.n1809 0.1295
R6114 VDD.n1108 VDD.n1107 0.1295
R6115 VDD.n1426 VDD.n1425 0.12875
R6116 VDD.n1103 VDD.n1102 0.128
R6117 VDD.n1919 VDD.n1918 0.128
R6118 VDD.n354 VDD.n353 0.128
R6119 VDD.n1923 VDD.n1922 0.128
R6120 VDD.n1999 VDD.n310 0.128
R6121 VDD.n2080 VDD.n2079 0.128
R6122 VDD.n2084 VDD.n2083 0.128
R6123 VDD.n772 VDD.n771 0.128
R6124 VDD.n2252 VDD.n2251 0.128
R6125 VDD.n180 VDD.n179 0.126816
R6126 VDD.n184 VDD.n183 0.126816
R6127 VDD.n1105 VDD.n1104 0.1265
R6128 VDD.n1682 VDD.n1681 0.12575
R6129 VDD.n1680 VDD.n1679 0.12575
R6130 VDD.n1828 VDD.n1827 0.12575
R6131 VDD.n1577 VDD.n498 0.125
R6132 VDD.n1740 VDD.n407 0.125
R6133 VDD.n1919 VDD.n320 0.125
R6134 VDD.n1922 VDD.n318 0.125
R6135 VDD.n2027 VDD.n2026 0.125
R6136 VDD.n2080 VDD.n253 0.125
R6137 VDD.n2083 VDD.n251 0.125
R6138 VDD.n773 VDD.n772 0.125
R6139 VDD.n2252 VDD.n222 0.125
R6140 VDD.n2255 VDD.n220 0.125
R6141 VDD.n49 VDD.n48 0.124975
R6142 VDD.n61 VDD.n60 0.124975
R6143 VDD.n73 VDD.n72 0.124975
R6144 VDD.n85 VDD.n84 0.124975
R6145 VDD.n97 VDD.n96 0.124975
R6146 VDD.n2051 VDD.n2050 0.12425
R6147 VDD.n2036 VDD.n2035 0.12425
R6148 VDD.n2168 VDD.n2167 0.12425
R6149 VDD.n152 VDD.n139 0.12425
R6150 VDD.n1834 VDD.n1833 0.1235
R6151 VDD.n542 VDD.n541 0.122
R6152 VDD.n1764 VDD.n1763 0.1205
R6153 VDD.n1766 VDD.n1765 0.1205
R6154 VDD.n1887 VDD.n1886 0.1205
R6155 VDD.n1453 VDD.n1452 0.119
R6156 VDD.n1301 VDD.n1300 0.119
R6157 VDD.n1664 VDD.n1663 0.1175
R6158 VDD.n1994 VDD.n1993 0.1175
R6159 VDD.n1564 VDD.n1563 0.11675
R6160 VDD.n1550 VDD.n1549 0.11675
R6161 VDD.n1179 VDD.n1178 0.11675
R6162 VDD.n2134 VDD.n2133 0.11675
R6163 VDD.n2133 VDD.n2132 0.116
R6164 VDD.n1460 VDD.n1459 0.1145
R6165 VDD.n1475 VDD.n1474 0.1145
R6166 VDD.n1330 VDD.n1329 0.1145
R6167 VDD.n1245 VDD.n1244 0.1145
R6168 VDD.n1227 VDD.n1226 0.1145
R6169 VDD.n1709 VDD.n1708 0.1145
R6170 VDD.n1204 VDD.n1203 0.1145
R6171 VDD.n1774 VDD.n1767 0.1145
R6172 VDD.n1158 VDD.n1157 0.1145
R6173 VDD.n1140 VDD.n1139 0.1145
R6174 VDD.n1072 VDD.n1071 0.1145
R6175 VDD.n1054 VDD.n1053 0.1145
R6176 VDD.n1914 VDD.n1913 0.1145
R6177 VDD.n1910 VDD.n1909 0.1145
R6178 VDD.n1025 VDD.n1024 0.1145
R6179 VDD.n1007 VDD.n1006 0.1145
R6180 VDD.n1928 VDD.n1927 0.1145
R6181 VDD.n978 VDD.n977 0.1145
R6182 VDD.n960 VDD.n959 0.1145
R6183 VDD.n898 VDD.n897 0.1145
R6184 VDD.n880 VDD.n879 0.1145
R6185 VDD.n2075 VDD.n2074 0.1145
R6186 VDD.n851 VDD.n850 0.1145
R6187 VDD.n833 VDD.n832 0.1145
R6188 VDD.n2089 VDD.n2088 0.1145
R6189 VDD.n804 VDD.n803 0.1145
R6190 VDD.n786 VDD.n785 0.1145
R6191 VDD.n767 VDD.n766 0.1145
R6192 VDD.n749 VDD.n748 0.1145
R6193 VDD.n725 VDD.n724 0.1145
R6194 VDD.n707 VDD.n706 0.1145
R6195 VDD.n2247 VDD.n2246 0.1145
R6196 VDD.n2229 VDD.n2228 0.1145
R6197 VDD.n2210 VDD.n2209 0.1145
R6198 VDD.n2194 VDD.n2193 0.1145
R6199 VDD.n545 VDD.n544 0.11375
R6200 VDD.n1908 VDD.n1907 0.11375
R6201 VDD.n1538 VDD.n1537 0.11225
R6202 VDD.n923 VDD.n307 0.11225
R6203 VDD.n1506 VDD.n548 0.1115
R6204 VDD.n109 VDD.n1 0.111156
R6205 VDD.n1438 VDD.n1437 0.10925
R6206 VDD.n2144 VDD.n2143 0.10925
R6207 VDD.n1423 VDD.n1422 0.1085
R6208 VDD.n1435 VDD.n1434 0.1085
R6209 VDD.n1472 VDD.n1471 0.1085
R6210 VDD.n1478 VDD.n1477 0.1085
R6211 VDD.n1496 VDD.n1495 0.1085
R6212 VDD.n1398 VDD.n500 0.1085
R6213 VDD.n1573 VDD.n1572 0.1085
R6214 VDD.n1532 VDD.n1531 0.1085
R6215 VDD.n1366 VDD.n1365 0.1085
R6216 VDD.n1594 VDD.n1593 0.1085
R6217 VDD.n1623 VDD.n1622 0.1085
R6218 VDD.n1278 VDD.n1277 0.1085
R6219 VDD.n1647 VDD.n1646 0.1085
R6220 VDD.n1727 VDD.n1726 0.1085
R6221 VDD.n1687 VDD.n1686 0.1085
R6222 VDD.n1826 VDD.n1825 0.1085
R6223 VDD.n1806 VDD.n1805 0.1085
R6224 VDD.n1101 VDD.n378 0.1085
R6225 VDD.n1853 VDD.n1852 0.1085
R6226 VDD.n1876 VDD.n1875 0.1085
R6227 VDD.n352 VDD.n351 0.1085
R6228 VDD.n1946 VDD.n1945 0.1085
R6229 VDD.n1997 VDD.n1996 0.1085
R6230 VDD.n2014 VDD.n2013 0.1085
R6231 VDD.n2056 VDD.n2055 0.1085
R6232 VDD.n2053 VDD.n2052 0.1085
R6233 VDD.n2037 VDD.n2036 0.1085
R6234 VDD.n2130 VDD.n2129 0.1085
R6235 VDD.n1649 VDD.n1648 0.10775
R6236 VDD.n1715 VDD.n1714 0.10775
R6237 VDD.n1371 VDD.n1370 0.107
R6238 VDD.n187 VDD.n175 0.10684
R6239 VDD.n12 VDD.n11 0.105754
R6240 VDD.n25 VDD.n24 0.105754
R6241 VDD.n37 VDD.n36 0.105754
R6242 VDD.n48 VDD.n47 0.105754
R6243 VDD.n60 VDD.n59 0.105754
R6244 VDD.n72 VDD.n71 0.105754
R6245 VDD.n84 VDD.n83 0.105754
R6246 VDD.n96 VDD.n95 0.105754
R6247 VDD.n1553 VDD.n1552 0.1055
R6248 VDD.n1574 VDD.n500 0.10475
R6249 VDD.n1714 VDD.n1713 0.10475
R6250 VDD.n1712 VDD.n1711 0.10475
R6251 VDD.n1111 VDD.n1110 0.1025
R6252 VDD.n1847 VDD.n1846 0.1025
R6253 VDD.n1883 VDD.n1882 0.10025
R6254 VDD.n633 VDD.n632 0.0995
R6255 VDD.n1445 VDD.n1444 0.0995
R6256 VDD.n1832 VDD.n1831 0.0995
R6257 VDD.n1498 VDD.n1497 0.09875
R6258 VDD.n1904 VDD.n1903 0.09875
R6259 VDD.n185 VDD.n184 0.0983947
R6260 VDD.n11 VDD.n10 0.0981271
R6261 VDD.n10 VDD.n9 0.0981271
R6262 VDD.n9 VDD.n8 0.0981271
R6263 VDD.n24 VDD.n23 0.0981271
R6264 VDD.n23 VDD.n22 0.0981271
R6265 VDD.n22 VDD.n21 0.0981271
R6266 VDD.n36 VDD.n35 0.0981271
R6267 VDD.n35 VDD.n34 0.0981271
R6268 VDD.n34 VDD.n33 0.0981271
R6269 VDD.n47 VDD.n46 0.0981271
R6270 VDD.n46 VDD.n45 0.0981271
R6271 VDD.n45 VDD.n44 0.0981271
R6272 VDD.n59 VDD.n58 0.0981271
R6273 VDD.n58 VDD.n57 0.0981271
R6274 VDD.n57 VDD.n56 0.0981271
R6275 VDD.n71 VDD.n70 0.0981271
R6276 VDD.n70 VDD.n69 0.0981271
R6277 VDD.n69 VDD.n68 0.0981271
R6278 VDD.n83 VDD.n82 0.0981271
R6279 VDD.n82 VDD.n81 0.0981271
R6280 VDD.n81 VDD.n80 0.0981271
R6281 VDD.n95 VDD.n94 0.0981271
R6282 VDD.n94 VDD.n93 0.0981271
R6283 VDD.n93 VDD.n92 0.0981271
R6284 VDD.n1533 VDD.n1532 0.098
R6285 VDD.n2043 VDD.n2042 0.098
R6286 VDD.n2149 VDD.n2148 0.098
R6287 VDD.n1589 VDD.n1588 0.0965
R6288 VDD.n1948 VDD.n1940 0.0965
R6289 VDD.n1473 VDD.n1472 0.09575
R6290 VDD.n1559 VDD.n1558 0.09425
R6291 VDD.n1978 VDD.n1977 0.09425
R6292 VDD.n290 VDD.n289 0.09425
R6293 VDD.n1510 VDD.n1509 0.0935
R6294 VDD.n1614 VDD.n1613 0.0935
R6295 VDD.n1297 VDD.n1296 0.0935
R6296 VDD.n1279 VDD.n1278 0.0935
R6297 VDD.n1726 VDD.n1725 0.0935
R6298 VDD.n1704 VDD.n1703 0.0935
R6299 VDD.n1702 VDD.n1701 0.0935
R6300 VDD.n1861 VDD.n1860 0.0935
R6301 VDD.n1968 VDD.n1967 0.0935
R6302 VDD.n2065 VDD.n2064 0.0935
R6303 VDD.n280 VDD.n279 0.0935
R6304 VDD.n2031 VDD.n293 0.09275
R6305 VDD.n1586 VDD.n1585 0.0905
R6306 VDD.n2123 VDD.n2122 0.0905
R6307 VDD.n1697 VDD.n1696 0.08975
R6308 VDD.n2017 VDD.n2016 0.08975
R6309 VDD.n119 VDD.n113 0.0896818
R6310 VDD.n1935 VDD.n1934 0.08825
R6311 VDD.n1982 VDD.n1981 0.08825
R6312 VDD.n1674 VDD.n1673 0.0875
R6313 VDD.n1289 VDD.n1288 0.08675
R6314 VDD.n1947 VDD.n1946 0.08675
R6315 VDD.n166 VDD.n135 0.08675
R6316 VDD.n2054 VDD.n2053 0.086
R6317 VDD.n2191 VDD.n229 0.086
R6318 VDD.n2301 VDD.n2300 0.086
R6319 VDD.n1310 VDD.n1309 0.08525
R6320 VDD.n1117 VDD.n1116 0.08525
R6321 VDD.n625 VDD.n624 0.0845
R6322 VDD.n627 VDD.n626 0.0845
R6323 VDD.n629 VDD.n628 0.0845
R6324 VDD.n631 VDD.n630 0.0845
R6325 VDD.n1447 VDD.n1446 0.0845
R6326 VDD.n1449 VDD.n1448 0.0845
R6327 VDD.n1451 VDD.n1450 0.0845
R6328 VDD.n1507 VDD.n1505 0.0845
R6329 VDD.n1378 VDD.n1377 0.0845
R6330 VDD.n1376 VDD.n1373 0.0845
R6331 VDD.n1261 VDD.n1260 0.0845
R6332 VDD.n1259 VDD.n1258 0.0845
R6333 VDD.n1257 VDD.n1256 0.0845
R6334 VDD.n1255 VDD.n1254 0.0845
R6335 VDD.n1253 VDD.n1252 0.0845
R6336 VDD.n1251 VDD.n1250 0.0845
R6337 VDD.n1249 VDD.n1248 0.0845
R6338 VDD.n1328 VDD.n1327 0.0845
R6339 VDD.n1326 VDD.n1325 0.0845
R6340 VDD.n1324 VDD.n1323 0.0845
R6341 VDD.n1322 VDD.n1321 0.0845
R6342 VDD.n1320 VDD.n1319 0.0845
R6343 VDD.n1318 VDD.n1317 0.0845
R6344 VDD.n1316 VDD.n1315 0.0845
R6345 VDD.n1314 VDD.n1313 0.0845
R6346 VDD.n1659 VDD.n1658 0.0845
R6347 VDD.n1220 VDD.n1219 0.0845
R6348 VDD.n1218 VDD.n1217 0.0845
R6349 VDD.n1216 VDD.n1215 0.0845
R6350 VDD.n1214 VDD.n1213 0.0845
R6351 VDD.n1212 VDD.n1211 0.0845
R6352 VDD.n1210 VDD.n1209 0.0845
R6353 VDD.n1208 VDD.n1207 0.0845
R6354 VDD.n1243 VDD.n1242 0.0845
R6355 VDD.n1241 VDD.n1240 0.0845
R6356 VDD.n1239 VDD.n1238 0.0845
R6357 VDD.n1237 VDD.n1236 0.0845
R6358 VDD.n1235 VDD.n1234 0.0845
R6359 VDD.n1233 VDD.n1232 0.0845
R6360 VDD.n1231 VDD.n1230 0.0845
R6361 VDD.n1229 VDD.n1228 0.0845
R6362 VDD.n1174 VDD.n1173 0.0845
R6363 VDD.n1172 VDD.n1171 0.0845
R6364 VDD.n1170 VDD.n1169 0.0845
R6365 VDD.n1168 VDD.n1167 0.0845
R6366 VDD.n1166 VDD.n1165 0.0845
R6367 VDD.n1164 VDD.n1163 0.0845
R6368 VDD.n1162 VDD.n1161 0.0845
R6369 VDD.n1772 VDD.n1771 0.0845
R6370 VDD.n1823 VDD.n1822 0.0845
R6371 VDD.n1821 VDD.n1820 0.0845
R6372 VDD.n1819 VDD.n1818 0.0845
R6373 VDD.n1817 VDD.n1816 0.0845
R6374 VDD.n1815 VDD.n1814 0.0845
R6375 VDD.n1813 VDD.n1812 0.0845
R6376 VDD.n1811 VDD.n1810 0.0845
R6377 VDD.n1088 VDD.n1087 0.0845
R6378 VDD.n1086 VDD.n1085 0.0845
R6379 VDD.n1084 VDD.n1083 0.0845
R6380 VDD.n1082 VDD.n1081 0.0845
R6381 VDD.n1080 VDD.n1079 0.0845
R6382 VDD.n1078 VDD.n1077 0.0845
R6383 VDD.n1076 VDD.n1075 0.0845
R6384 VDD.n1156 VDD.n1155 0.0845
R6385 VDD.n1154 VDD.n1153 0.0845
R6386 VDD.n1152 VDD.n1151 0.0845
R6387 VDD.n1150 VDD.n1149 0.0845
R6388 VDD.n1148 VDD.n1147 0.0845
R6389 VDD.n1146 VDD.n1145 0.0845
R6390 VDD.n1144 VDD.n1143 0.0845
R6391 VDD.n1142 VDD.n1141 0.0845
R6392 VDD.n1138 VDD.n1137 0.0845
R6393 VDD.n1136 VDD.n1135 0.0845
R6394 VDD.n1134 VDD.n1133 0.0845
R6395 VDD.n1132 VDD.n1131 0.0845
R6396 VDD.n1130 VDD.n1129 0.0845
R6397 VDD.n1128 VDD.n1127 0.0845
R6398 VDD.n1125 VDD.n1124 0.0845
R6399 VDD.n1123 VDD.n1122 0.0845
R6400 VDD.n1041 VDD.n1040 0.0845
R6401 VDD.n1039 VDD.n1038 0.0845
R6402 VDD.n1037 VDD.n1036 0.0845
R6403 VDD.n1035 VDD.n1034 0.0845
R6404 VDD.n1033 VDD.n1032 0.0845
R6405 VDD.n1031 VDD.n1030 0.0845
R6406 VDD.n1029 VDD.n1028 0.0845
R6407 VDD.n1070 VDD.n1069 0.0845
R6408 VDD.n1068 VDD.n1067 0.0845
R6409 VDD.n1066 VDD.n1065 0.0845
R6410 VDD.n1064 VDD.n1063 0.0845
R6411 VDD.n1062 VDD.n1061 0.0845
R6412 VDD.n1060 VDD.n1059 0.0845
R6413 VDD.n1058 VDD.n1057 0.0845
R6414 VDD.n1056 VDD.n1055 0.0845
R6415 VDD.n1052 VDD.n1051 0.0845
R6416 VDD.n1050 VDD.n1049 0.0845
R6417 VDD.n1048 VDD.n1047 0.0845
R6418 VDD.n1046 VDD.n1045 0.0845
R6419 VDD.n1044 VDD.n1043 0.0845
R6420 VDD.n1042 VDD.n320 0.0845
R6421 VDD.n1918 VDD.n1917 0.0845
R6422 VDD.n1916 VDD.n1915 0.0845
R6423 VDD.n994 VDD.n993 0.0845
R6424 VDD.n992 VDD.n991 0.0845
R6425 VDD.n990 VDD.n989 0.0845
R6426 VDD.n988 VDD.n987 0.0845
R6427 VDD.n986 VDD.n985 0.0845
R6428 VDD.n984 VDD.n983 0.0845
R6429 VDD.n982 VDD.n981 0.0845
R6430 VDD.n1023 VDD.n1022 0.0845
R6431 VDD.n1021 VDD.n1020 0.0845
R6432 VDD.n1019 VDD.n1018 0.0845
R6433 VDD.n1017 VDD.n1016 0.0845
R6434 VDD.n1015 VDD.n1014 0.0845
R6435 VDD.n1013 VDD.n1012 0.0845
R6436 VDD.n1011 VDD.n1010 0.0845
R6437 VDD.n1009 VDD.n1008 0.0845
R6438 VDD.n1005 VDD.n1004 0.0845
R6439 VDD.n1003 VDD.n1002 0.0845
R6440 VDD.n1001 VDD.n1000 0.0845
R6441 VDD.n999 VDD.n998 0.0845
R6442 VDD.n997 VDD.n996 0.0845
R6443 VDD.n995 VDD.n318 0.0845
R6444 VDD.n1924 VDD.n1923 0.0845
R6445 VDD.n1926 VDD.n1925 0.0845
R6446 VDD.n914 VDD.n913 0.0845
R6447 VDD.n912 VDD.n911 0.0845
R6448 VDD.n910 VDD.n909 0.0845
R6449 VDD.n908 VDD.n907 0.0845
R6450 VDD.n906 VDD.n905 0.0845
R6451 VDD.n904 VDD.n903 0.0845
R6452 VDD.n902 VDD.n901 0.0845
R6453 VDD.n976 VDD.n975 0.0845
R6454 VDD.n974 VDD.n973 0.0845
R6455 VDD.n972 VDD.n971 0.0845
R6456 VDD.n970 VDD.n969 0.0845
R6457 VDD.n968 VDD.n967 0.0845
R6458 VDD.n966 VDD.n965 0.0845
R6459 VDD.n964 VDD.n963 0.0845
R6460 VDD.n962 VDD.n961 0.0845
R6461 VDD.n958 VDD.n957 0.0845
R6462 VDD.n956 VDD.n955 0.0845
R6463 VDD.n954 VDD.n953 0.0845
R6464 VDD.n952 VDD.n951 0.0845
R6465 VDD.n950 VDD.n949 0.0845
R6466 VDD.n948 VDD.n947 0.0845
R6467 VDD.n945 VDD.n944 0.0845
R6468 VDD.n943 VDD.n942 0.0845
R6469 VDD.n940 VDD.n939 0.0845
R6470 VDD.n938 VDD.n937 0.0845
R6471 VDD.n936 VDD.n935 0.0845
R6472 VDD.n934 VDD.n933 0.0845
R6473 VDD.n867 VDD.n866 0.0845
R6474 VDD.n865 VDD.n864 0.0845
R6475 VDD.n863 VDD.n862 0.0845
R6476 VDD.n861 VDD.n860 0.0845
R6477 VDD.n859 VDD.n858 0.0845
R6478 VDD.n857 VDD.n856 0.0845
R6479 VDD.n855 VDD.n854 0.0845
R6480 VDD.n896 VDD.n895 0.0845
R6481 VDD.n894 VDD.n893 0.0845
R6482 VDD.n892 VDD.n891 0.0845
R6483 VDD.n890 VDD.n889 0.0845
R6484 VDD.n888 VDD.n887 0.0845
R6485 VDD.n886 VDD.n885 0.0845
R6486 VDD.n884 VDD.n883 0.0845
R6487 VDD.n882 VDD.n881 0.0845
R6488 VDD.n878 VDD.n877 0.0845
R6489 VDD.n876 VDD.n875 0.0845
R6490 VDD.n874 VDD.n873 0.0845
R6491 VDD.n872 VDD.n871 0.0845
R6492 VDD.n870 VDD.n869 0.0845
R6493 VDD.n868 VDD.n253 0.0845
R6494 VDD.n2079 VDD.n2078 0.0845
R6495 VDD.n2077 VDD.n2076 0.0845
R6496 VDD.n820 VDD.n819 0.0845
R6497 VDD.n818 VDD.n817 0.0845
R6498 VDD.n816 VDD.n815 0.0845
R6499 VDD.n814 VDD.n813 0.0845
R6500 VDD.n812 VDD.n811 0.0845
R6501 VDD.n810 VDD.n809 0.0845
R6502 VDD.n808 VDD.n807 0.0845
R6503 VDD.n849 VDD.n848 0.0845
R6504 VDD.n847 VDD.n846 0.0845
R6505 VDD.n845 VDD.n844 0.0845
R6506 VDD.n843 VDD.n842 0.0845
R6507 VDD.n841 VDD.n840 0.0845
R6508 VDD.n839 VDD.n838 0.0845
R6509 VDD.n837 VDD.n836 0.0845
R6510 VDD.n835 VDD.n834 0.0845
R6511 VDD.n831 VDD.n830 0.0845
R6512 VDD.n829 VDD.n828 0.0845
R6513 VDD.n827 VDD.n826 0.0845
R6514 VDD.n825 VDD.n824 0.0845
R6515 VDD.n823 VDD.n822 0.0845
R6516 VDD.n821 VDD.n251 0.0845
R6517 VDD.n2085 VDD.n2084 0.0845
R6518 VDD.n2087 VDD.n2086 0.0845
R6519 VDD.n741 VDD.n740 0.0845
R6520 VDD.n739 VDD.n738 0.0845
R6521 VDD.n737 VDD.n736 0.0845
R6522 VDD.n735 VDD.n734 0.0845
R6523 VDD.n733 VDD.n732 0.0845
R6524 VDD.n731 VDD.n730 0.0845
R6525 VDD.n729 VDD.n728 0.0845
R6526 VDD.n802 VDD.n801 0.0845
R6527 VDD.n800 VDD.n799 0.0845
R6528 VDD.n798 VDD.n797 0.0845
R6529 VDD.n796 VDD.n795 0.0845
R6530 VDD.n794 VDD.n793 0.0845
R6531 VDD.n792 VDD.n791 0.0845
R6532 VDD.n790 VDD.n789 0.0845
R6533 VDD.n788 VDD.n787 0.0845
R6534 VDD.n784 VDD.n783 0.0845
R6535 VDD.n782 VDD.n781 0.0845
R6536 VDD.n780 VDD.n779 0.0845
R6537 VDD.n778 VDD.n777 0.0845
R6538 VDD.n776 VDD.n775 0.0845
R6539 VDD.n774 VDD.n773 0.0845
R6540 VDD.n771 VDD.n770 0.0845
R6541 VDD.n769 VDD.n768 0.0845
R6542 VDD.n765 VDD.n764 0.0845
R6543 VDD.n763 VDD.n762 0.0845
R6544 VDD.n761 VDD.n760 0.0845
R6545 VDD.n759 VDD.n758 0.0845
R6546 VDD.n757 VDD.n756 0.0845
R6547 VDD.n755 VDD.n754 0.0845
R6548 VDD.n753 VDD.n752 0.0845
R6549 VDD.n751 VDD.n750 0.0845
R6550 VDD.n747 VDD.n746 0.0845
R6551 VDD.n745 VDD.n744 0.0845
R6552 VDD.n743 VDD.n742 0.0845
R6553 VDD.n2155 VDD.n2154 0.0845
R6554 VDD.n2157 VDD.n2156 0.0845
R6555 VDD.n2163 VDD.n2162 0.0845
R6556 VDD.n694 VDD.n693 0.0845
R6557 VDD.n692 VDD.n691 0.0845
R6558 VDD.n690 VDD.n689 0.0845
R6559 VDD.n688 VDD.n687 0.0845
R6560 VDD.n686 VDD.n685 0.0845
R6561 VDD.n684 VDD.n683 0.0845
R6562 VDD.n682 VDD.n681 0.0845
R6563 VDD.n723 VDD.n722 0.0845
R6564 VDD.n721 VDD.n720 0.0845
R6565 VDD.n719 VDD.n718 0.0845
R6566 VDD.n717 VDD.n716 0.0845
R6567 VDD.n715 VDD.n714 0.0845
R6568 VDD.n713 VDD.n712 0.0845
R6569 VDD.n711 VDD.n710 0.0845
R6570 VDD.n709 VDD.n708 0.0845
R6571 VDD.n705 VDD.n704 0.0845
R6572 VDD.n703 VDD.n702 0.0845
R6573 VDD.n701 VDD.n700 0.0845
R6574 VDD.n699 VDD.n698 0.0845
R6575 VDD.n697 VDD.n696 0.0845
R6576 VDD.n695 VDD.n222 0.0845
R6577 VDD.n2251 VDD.n2250 0.0845
R6578 VDD.n2249 VDD.n2248 0.0845
R6579 VDD.n2245 VDD.n2244 0.0845
R6580 VDD.n2243 VDD.n2242 0.0845
R6581 VDD.n2241 VDD.n2240 0.0845
R6582 VDD.n2239 VDD.n2238 0.0845
R6583 VDD.n2237 VDD.n2236 0.0845
R6584 VDD.n2235 VDD.n2234 0.0845
R6585 VDD.n2233 VDD.n2232 0.0845
R6586 VDD.n2231 VDD.n2230 0.0845
R6587 VDD.n2227 VDD.n2226 0.0845
R6588 VDD.n2225 VDD.n2224 0.0845
R6589 VDD.n2223 VDD.n2222 0.0845
R6590 VDD.n2221 VDD.n2220 0.0845
R6591 VDD.n2218 VDD.n2217 0.0845
R6592 VDD.n2216 VDD.n2215 0.0845
R6593 VDD.n2214 VDD.n2213 0.0845
R6594 VDD.n2212 VDD.n2211 0.0845
R6595 VDD.n2198 VDD.n2197 0.0845
R6596 VDD.n2196 VDD.n2195 0.0845
R6597 VDD.n2318 VDD.n2317 0.0845
R6598 VDD.n108 VDD.n12 0.0843983
R6599 VDD.n26 VDD.n25 0.0843983
R6600 VDD.n1574 VDD.n1573 0.08375
R6601 VDD.n1528 VDD.n1527 0.08375
R6602 VDD.n2188 VDD.n231 0.083
R6603 VDD.n2302 VDD.n2301 0.083
R6604 VDD.n1717 VDD.n1716 0.08225
R6605 VDD.n1432 VDD.n1431 0.0815
R6606 VDD.n1749 VDD.n1748 0.0815
R6607 VDD.n1893 VDD.n1892 0.0815
R6608 VDD.n1888 VDD.n1887 0.0815
R6609 VDD.n1416 VDD.n1415 0.08075
R6610 VDD.n1595 VDD.n1594 0.08075
R6611 VDD.n1287 VDD.n1286 0.08075
R6612 VDD.n1691 VDD.n1690 0.08075
R6613 VDD.n2142 VDD.n2141 0.07925
R6614 VDD.n1700 VDD.n1699 0.0785
R6615 VDD.n1799 VDD.n1798 0.0785
R6616 VDD.n1355 VDD.n1354 0.07775
R6617 VDD.n1544 VDD.n1543 0.077
R6618 VDD.n98 VDD.n26 0.0755336
R6619 VDD.n1464 VDD.n1463 0.0755
R6620 VDD.n540 VDD.n539 0.0755
R6621 VDD.n1842 VDD.n1841 0.0755
R6622 VDD.n1859 VDD.n1858 0.0755
R6623 VDD.n2022 VDD.n2021 0.07475
R6624 VDD.n1568 VDD.n1567 0.0725
R6625 VDD.n1767 VDD.n1766 0.0725
R6626 VDD.n1523 VDD.n1522 0.071
R6627 VDD.n1639 VDD.n1638 0.071
R6628 VDD.n1881 VDD.n1880 0.07025
R6629 VDD.n2030 VDD.n2029 0.07025
R6630 VDD.n1454 VDD.n1453 0.0695
R6631 VDD.n1456 VDD.n1455 0.0695
R6632 VDD.n1492 VDD.n1491 0.0695
R6633 VDD.n1745 VDD.n1744 0.0695
R6634 VDD.n1747 VDD.n1746 0.0695
R6635 VDD.n2126 VDD.n2125 0.0695
R6636 VDD.n927 VDD.n926 0.068
R6637 VDD.n1503 VDD.n1502 0.06725
R6638 VDD.n1693 VDD.n1692 0.06575
R6639 VDD.n2139 VDD.n2138 0.065
R6640 VDD.n2125 VDD.n2124 0.065
R6641 VDD.n2153 VDD.n2152 0.065
R6642 VDD.n1441 VDD.n1440 0.06425
R6643 VDD.n1406 VDD.n1405 0.0635
R6644 VDD.n1750 VDD.n1749 0.06275
R6645 VDD.n679 VDD.n637 0.062
R6646 VDD.n1636 VDD.n1635 0.06125
R6647 VDD.n1277 VDD.n1276 0.0605
R6648 VDD.n1728 VDD.n1727 0.0605
R6649 VDD.n2120 VDD.n2119 0.0605
R6650 VDD.n101 VDD.n100 0.0595164
R6651 VDD.n102 VDD.n101 0.0595164
R6652 VDD.n102 VDD.n13 0.0595164
R6653 VDD.n106 VDD.n13 0.0595164
R6654 VDD.n107 VDD.n106 0.0595164
R6655 VDD.n1415 VDD.n1414 0.05825
R6656 VDD.n108 VDD.n107 0.0578934
R6657 VDD.n1430 VDD.n1429 0.0575
R6658 VDD.n1897 VDD.n1896 0.0575
R6659 VDD.n1584 VDD.n1583 0.05675
R6660 VDD.n1484 VDD.n1483 0.056
R6661 VDD.n1743 VDD.n405 0.056
R6662 VDD.n1308 VDD.n1307 0.05525
R6663 VDD.n1312 VDD.n1311 0.0545
R6664 VDD.n1121 VDD.n1120 0.0545
R6665 VDD.n1992 VDD.n1991 0.0545
R6666 VDD.n941 VDD.n940 0.0545
R6667 VDD.n2015 VDD.n2014 0.0545
R6668 VDD.n2161 VDD.n2160 0.0545
R6669 VDD.n2173 VDD.n2172 0.0545
R6670 VDD.n1535 VDD.n1534 0.053
R6671 VDD.n1380 VDD.n1379 0.05225
R6672 VDD.n1466 VDD.n1465 0.0515
R6673 VDD.n1477 VDD.n1476 0.05075
R6674 VDD.n1495 VDD.n1494 0.05075
R6675 VDD.n1501 VDD.n1500 0.05075
R6676 VDD.n1298 VDD.n1297 0.05075
R6677 VDD.n1825 VDD.n1824 0.05075
R6678 VDD.n1711 VDD.n1710 0.05
R6679 VDD.n1695 VDD.n1694 0.05
R6680 VDD.n1940 VDD.n1939 0.05
R6681 VDD.n1561 VDD.n1560 0.04925
R6682 VDD.n1655 VDD.n1654 0.04925
R6683 VDD.n1667 VDD.n458 0.0485
R6684 VDD.n2020 VDD.n293 0.0485
R6685 VDD.n1752 VDD.n1751 0.04775
R6686 VDD.n1652 VDD.n1651 0.0455
R6687 VDD.n1641 VDD.n482 0.044
R6688 VDD.n2002 VDD.n307 0.044
R6689 VDD.n1855 VDD.n361 0.04325
R6690 VDD.n100 VDD.n26 0.0431393
R6691 VDD.n1284 VDD.n1283 0.0425
R6692 VDD.n119 VDD.n118 0.0422273
R6693 VDD.n1127 VDD.n1126 0.041
R6694 VDD.n947 VDD.n946 0.041
R6695 VDD.n1424 VDD.n1423 0.04025
R6696 VDD.n1551 VDD.n1550 0.04025
R6697 VDD.n1303 VDD.n1302 0.04025
R6698 VDD.n1838 VDD.n378 0.04025
R6699 VDD.n2062 VDD.n2061 0.04025
R6700 VDD.n635 VDD.n213 0.0396304
R6701 VDD.n2335 VDD.n2334 0.0396304
R6702 VDD.n1721 VDD.n1720 0.0395
R6703 VDD.n2007 VDD.n2006 0.0395
R6704 VDD.n1275 VDD.n479 0.038
R6705 VDD.n1844 VDD.n1843 0.0365
R6706 VDD.n2022 VDD.n2018 0.03425
R6707 VDD.n2136 VDD.n2135 0.03425
R6708 VDD.n1739 VDD.n1738 0.0335
R6709 VDD.n1737 VDD.n1736 0.0335
R6710 VDD.n1733 VDD.n1732 0.0335
R6711 VDD.n1723 VDD.n1722 0.0335
R6712 VDD.n1868 VDD.n1867 0.0335
R6713 VDD.n1975 VDD.n1974 0.0335
R6714 VDD.n287 VDD.n286 0.0335
R6715 VDD.n99 VDD.n14 0.0332273
R6716 VDD.n103 VDD.n14 0.0332273
R6717 VDD.n104 VDD.n103 0.0332273
R6718 VDD.n105 VDD.n104 0.0332273
R6719 VDD.n105 VDD.n1 0.0332273
R6720 VDD.n1411 VDD.n1410 0.03275
R6721 VDD.n1359 VDD.n1358 0.03275
R6722 VDD.n1540 VDD.n1539 0.0305
R6723 VDD.n1370 VDD.n1369 0.0305
R6724 VDD.n2102 VDD.n2098 0.0305
R6725 VDD.n676 VDD.n675 0.0305
R6726 VDD.n2259 VDD.n2258 0.0305
R6727 VDD.n2276 VDD.n2270 0.0305
R6728 VDD.n2320 VDD.n2319 0.0305
R6729 VDD.n1439 VDD.n1438 0.02975
R6730 VDD.n198 VDD.n124 0.0296828
R6731 VDD.n185 VDD.n180 0.0289211
R6732 VDD.n1115 VDD.n1114 0.02825
R6733 VDD.n1113 VDD.n1112 0.0275
R6734 VDD.n1890 VDD.n1889 0.0275
R6735 VDD.n2146 VDD.n2145 0.0275
R6736 VDD.n211 VDD.n121 0.0270738
R6737 VDD.n207 VDD.n121 0.0270738
R6738 VDD.n207 VDD.n206 0.0270738
R6739 VDD.n206 VDD.n205 0.0270738
R6740 VDD.n205 VDD.n123 0.0270738
R6741 VDD.n201 VDD.n123 0.0270738
R6742 VDD.n201 VDD.n200 0.0270738
R6743 VDD.n199 VDD.n125 0.0270738
R6744 VDD.n195 VDD.n125 0.0270738
R6745 VDD.n195 VDD.n194 0.0270738
R6746 VDD.n194 VDD.n193 0.0270738
R6747 VDD.n193 VDD.n127 0.0270738
R6748 VDD.n189 VDD.n127 0.0270738
R6749 VDD.n189 VDD.n188 0.0270738
R6750 VDD.n1306 VDD.n1305 0.02675
R6751 VDD.n1181 VDD.n1180 0.02675
R6752 VDD.n1459 VDD.n1458 0.0245
R6753 VDD.n1542 VDD.n1541 0.0245
R6754 VDD.n2315 VDD.n2314 0.0245
R6755 VDD.n1527 VDD.n1526 0.02375
R6756 VDD.n538 VDD.n537 0.023
R6757 VDD.n1580 VDD.n1579 0.023
R6758 VDD.n1331 VDD.n1330 0.023
R6759 VDD.n1246 VDD.n1245 0.023
R6760 VDD.n1205 VDD.n1204 0.023
R6761 VDD.n1159 VDD.n1158 0.023
R6762 VDD.n1073 VDD.n1072 0.023
R6763 VDD.n1026 VDD.n1025 0.023
R6764 VDD.n979 VDD.n978 0.023
R6765 VDD.n899 VDD.n898 0.023
R6766 VDD.n2035 VDD.n2034 0.023
R6767 VDD.n852 VDD.n851 0.023
R6768 VDD.n805 VDD.n804 0.023
R6769 VDD.n726 VDD.n725 0.023
R6770 VDD.n1290 VDD.n1289 0.0215
R6771 VDD.n1936 VDD.n1935 0.02075
R6772 VDD.n1981 VDD.n1980 0.02075
R6773 VDD.n1645 VDD.n1644 0.02
R6774 VDD.n2152 VDD.n239 0.02
R6775 VDD.n2220 VDD.n2219 0.02
R6776 VDD.n2331 VDD.n217 0.02
R6777 VDD.n1863 VDD.n1862 0.0185
R6778 VDD.n1970 VDD.n1969 0.0185
R6779 VDD.n282 VDD.n281 0.0185
R6780 VDD.n2046 VDD.n2045 0.017
R6781 VDD.n1296 VDD.n1295 0.0155
R6782 VDD.n1294 VDD.n1293 0.0155
R6783 VDD.n1668 VDD.n1665 0.01475
R6784 VDD.n187 VDD.n186 0.0143449
R6785 VDD.n212 VDD.n120 0.0142641
R6786 VDD.n451 VDD.n450 0.014
R6787 VDD.n1896 VDD.n1895 0.01325
R6788 VDD.n175 VDD.n129 0.0127117
R6789 VDD.n171 VDD.n129 0.0127117
R6790 VDD.n171 VDD.n170 0.0127117
R6791 VDD.n170 VDD.n169 0.0127117
R6792 VDD.n169 VDD.n131 0.0127117
R6793 VDD.n165 VDD.n131 0.0127117
R6794 VDD.n165 VDD.n164 0.0127117
R6795 VDD.n164 VDD.n136 0.0127117
R6796 VDD.n160 VDD.n136 0.0127117
R6797 VDD.n160 VDD.n159 0.0127117
R6798 VDD.n159 VDD.n158 0.0127117
R6799 VDD.n158 VDD.n138 0.0127117
R6800 VDD.n154 VDD.n138 0.0127117
R6801 VDD.n154 VDD.n153 0.0127117
R6802 VDD.n153 VDD.n140 0.0127117
R6803 VDD.n149 VDD.n140 0.0127117
R6804 VDD.n149 VDD.n148 0.0127117
R6805 VDD.n148 VDD.n147 0.0127117
R6806 VDD.n147 VDD.n0 0.0127117
R6807 VDD.n1106 VDD.n1105 0.0125
R6808 VDD.n1399 VDD.n1398 0.011
R6809 VDD.n1572 VDD.n1571 0.011
R6810 VDD.n930 VDD.n929 0.011
R6811 VDD.n1678 VDD.n1677 0.01025
R6812 VDD.n1856 VDD.n1853 0.01025
R6813 VDD.n623 VDD.n622 0.0095
R6814 VDD.n634 VDD.n633 0.0095
R6815 VDD.n1866 VDD.n1865 0.0095
R6816 VDD.n1973 VDD.n1972 0.0095
R6817 VDD.n285 VDD.n284 0.0095
R6818 VDD.n1364 VDD.n1363 0.008
R6819 VDD.n1835 VDD.n1834 0.008
R6820 VDD.n1805 VDD.n1804 0.0065
R6821 VDD.n1875 VDD.n1874 0.0065
R6822 VDD.n1688 VDD.n1687 0.00575
R6823 VDD.n1885 VDD.n1884 0.00575
R6824 VDD.n210 VDD.n209 0.00363095
R6825 VDD.n209 VDD.n208 0.00363095
R6826 VDD.n208 VDD.n122 0.00363095
R6827 VDD.n204 VDD.n122 0.00363095
R6828 VDD.n204 VDD.n203 0.00363095
R6829 VDD.n203 VDD.n202 0.00363095
R6830 VDD.n202 VDD.n124 0.00363095
R6831 VDD.n198 VDD.n197 0.00363095
R6832 VDD.n197 VDD.n196 0.00363095
R6833 VDD.n196 VDD.n126 0.00363095
R6834 VDD.n192 VDD.n126 0.00363095
R6835 VDD.n192 VDD.n191 0.00363095
R6836 VDD.n191 VDD.n190 0.00363095
R6837 VDD.n190 VDD.n128 0.00363095
R6838 VDD.n1403 VDD.n1402 0.0035
R6839 VDD.n1681 VDD.n1680 0.0035
R6840 VDD.n1735 VDD.n1734 0.0035
R6841 VDD.n1622 VDD.n1621 0.00275
R6842 VDD.n1901 VDD.n1900 0.00275
R6843 VDD.n210 VDD.n120 0.00206547
R6844 VDD.n186 VDD.n128 0.00206547
R6845 VDD.n1989 VDD.n1988 0.002
R6846 VDD.n1987 VDD.n1986 0.002
R6847 VSS.n2442 VSS.n2441 815620
R6848 VSS.n2441 VSS.n2440 386085
R6849 VSS.n2444 VSS.n2443 20110.8
R6850 VSS.n2446 VSS.n2445 20110.8
R6851 VSS.n2448 VSS.n2447 20110.8
R6852 VSS.n2450 VSS.n2449 20110.8
R6853 VSS.n2452 VSS.n2451 20110.8
R6854 VSS.n2454 VSS.n2453 20110.8
R6855 VSS.n2456 VSS.n2455 13165.9
R6856 VSS.n2534 VSS.t2083 8049.82
R6857 VSS.n2494 VSS.n30 6725.25
R6858 VSS.n2537 VSS.n2513 3732.14
R6859 VSS.n2534 VSS.n2516 3632.35
R6860 VSS.n2539 VSS.n2538 3421.91
R6861 VSS.n542 VSS.n30 3273.43
R6862 VSS.n30 VSS.n11 3166.67
R6863 VSS.n2536 VSS.n2514 2972.65
R6864 VSS.n2423 VSS.n2422 2580.82
R6865 VSS.t2252 VSS.t4290 2506.75
R6866 VSS.t1483 VSS.t4191 2419.03
R6867 VSS.n578 VSS.n542 2318.66
R6868 VSS.n2232 VSS.n2231 2175.84
R6869 VSS.n2218 VSS.n2217 2138.68
R6870 VSS.t4048 VSS.t1629 2105.11
R6871 VSS.t2716 VSS.n369 2086.65
R6872 VSS.n2535 VSS.n2515 2077.22
R6873 VSS.t4095 VSS.t2637 2068.18
R6874 VSS.t2637 VSS.t3289 2068.18
R6875 VSS.t3289 VSS.t1942 2068.18
R6876 VSS.t1942 VSS.t2556 2068.18
R6877 VSS.t2556 VSS.t3012 2068.18
R6878 VSS.t3012 VSS.t1287 2068.18
R6879 VSS.t1287 VSS.t2193 2068.18
R6880 VSS.t2193 VSS.t1164 2068.18
R6881 VSS.t2353 VSS.t4024 2068.18
R6882 VSS.t2184 VSS.t1089 2068.18
R6883 VSS.t1489 VSS.t2184 2068.18
R6884 VSS.t367 VSS.t541 2068.18
R6885 VSS.t3629 VSS.t2260 2068.18
R6886 VSS.t3629 VSS.t1668 2068.18
R6887 VSS.t2137 VSS.t2597 2068.18
R6888 VSS.t3040 VSS.t1871 2068.18
R6889 VSS.t1871 VSS.t3022 2068.18
R6890 VSS.t3022 VSS.t4126 2068.18
R6891 VSS.t4126 VSS.t1745 2068.18
R6892 VSS.t2120 VSS.t4212 2068.18
R6893 VSS.t4212 VSS.t2855 2068.18
R6894 VSS.t2855 VSS.t2248 2068.18
R6895 VSS.t2248 VSS.t1491 2068.18
R6896 VSS.t1491 VSS.t1475 2068.18
R6897 VSS.t1475 VSS.t2256 2068.18
R6898 VSS.t2256 VSS.t4153 2068.18
R6899 VSS.t4153 VSS.t2831 2068.18
R6900 VSS.t529 VSS.t477 2068.18
R6901 VSS.t1883 VSS.t967 2068.18
R6902 VSS.t3730 VSS.t1425 2068.18
R6903 VSS.t4255 VSS.t2779 2068.18
R6904 VSS.t3918 VSS.t665 2068.18
R6905 VSS.t1566 VSS.t2191 2068.18
R6906 VSS.t1511 VSS.t4108 2068.18
R6907 VSS.t2213 VSS.t2653 2068.18
R6908 VSS.t1141 VSS.t2716 2068.18
R6909 VSS.t2231 VSS.t1141 2068.18
R6910 VSS.t1265 VSS.t2231 2068.18
R6911 VSS.t1270 VSS.t1265 2068.18
R6912 VSS.t1559 VSS.t1270 2068.18
R6913 VSS.t3293 VSS.t1559 2068.18
R6914 VSS.t1768 VSS.t3504 2068.18
R6915 VSS.t3504 VSS.t2400 2068.18
R6916 VSS.t2400 VSS.t3856 2068.18
R6917 VSS.n2126 VSS.t2500 2064.13
R6918 VSS.t2220 VSS.t901 1925.07
R6919 VSS.n2133 VSS.t1312 1901.99
R6920 VSS.t1242 VSS.t825 1883.52
R6921 VSS.n1716 VSS.t695 1883.52
R6922 VSS.t532 VSS.t2065 1883.52
R6923 VSS.t795 VSS.t3239 1883.52
R6924 VSS.t1899 VSS.t1210 1883.52
R6925 VSS.t3856 VSS.t3878 1883.52
R6926 VSS.t676 VSS.t2599 1846.59
R6927 VSS.t4184 VSS.t2318 1809.66
R6928 VSS.t3682 VSS.t508 1805.04
R6929 VSS.t4299 VSS.t3330 1805.04
R6930 VSS.t3838 VSS.t360 1781.96
R6931 VSS.t3295 VSS.t4316 1768.11
R6932 VSS.n2538 VSS.n11 1761.11
R6933 VSS.t3858 VSS.t3104 1758.88
R6934 VSS.t313 VSS.n71 1754.26
R6935 VSS.n579 VSS.t555 1754.26
R6936 VSS.t2522 VSS.t516 1754.26
R6937 VSS.t2355 VSS.t9 1735.8
R6938 VSS.t3670 VSS.t4136 1735.8
R6939 VSS.n2125 VSS.t852 1735.8
R6940 VSS.t3908 VSS.t1155 1735.8
R6941 VSS.t686 VSS.t3944 1731.18
R6942 VSS.t3637 VSS.t836 1731.18
R6943 VSS.t1322 VSS.t2930 1717.33
R6944 VSS.t969 VSS.t1555 1717.33
R6945 VSS.t1854 VSS.t1525 1717.33
R6946 VSS.t2517 VSS.t1642 1717.33
R6947 VSS.n2536 VSS.n2535 1712.04
R6948 VSS.t2169 VSS.t486 1698.86
R6949 VSS.t4142 VSS.t4225 1698.86
R6950 VSS.t3373 VSS.t10 1698.86
R6951 VSS.t4204 VSS.t1934 1698.86
R6952 VSS.t4208 VSS.t3310 1698.86
R6953 VSS.t370 VSS.t4190 1698.86
R6954 VSS.t2309 VSS.t2520 1685.01
R6955 VSS.t3381 VSS.t4116 1638.85
R6956 VSS.n2535 VSS.n2534 1635.19
R6957 VSS.n2424 VSS.n2423 1626
R6958 VSS.t903 VSS.t1994 1620.38
R6959 VSS.t1196 VSS.t2414 1620.38
R6960 VSS.t3051 VSS.t3680 1620.38
R6961 VSS.t4135 VSS.t3589 1588.07
R6962 VSS.t2020 VSS.t2918 1588.07
R6963 VSS.t1024 VSS.t1016 1588.07
R6964 VSS.n94 VSS.t2927 1569.6
R6965 VSS.t1164 VSS.n76 1569.6
R6966 VSS.t3486 VSS.n359 1569.6
R6967 VSS.t3057 VSS.n75 1569.6
R6968 VSS.t2081 VSS.n360 1569.6
R6969 VSS.t1745 VSS.n74 1569.6
R6970 VSS.t3125 VSS.n361 1569.6
R6971 VSS.t2055 VSS.n73 1569.6
R6972 VSS.t3502 VSS.n362 1569.6
R6973 VSS.t3059 VSS.n363 1569.6
R6974 VSS.t3397 VSS.n364 1569.6
R6975 VSS.t2592 VSS.n365 1569.6
R6976 VSS.t4353 VSS.n366 1569.6
R6977 VSS.t1891 VSS.n367 1569.6
R6978 VSS.t4357 VSS.n368 1569.6
R6979 VSS.t2312 VSS.n370 1569.6
R6980 VSS.t2096 VSS.n371 1569.6
R6981 VSS.n2438 VSS.n2437 1566.07
R6982 VSS.n2435 VSS.n2434 1566.07
R6983 VSS.n2430 VSS.n2429 1566.07
R6984 VSS.n2427 VSS.n2426 1566.07
R6985 VSS.t3888 VSS.t3904 1551.14
R6986 VSS.t977 VSS.t1973 1551.14
R6987 VSS.t1698 VSS.t3036 1551.14
R6988 VSS.t3476 VSS.t3147 1551.14
R6989 VSS.t2651 VSS.t2884 1551.14
R6990 VSS.t3970 VSS.t4001 1551.14
R6991 VSS.t3933 VSS.t2454 1551.14
R6992 VSS.t3974 VSS.t3933 1551.14
R6993 VSS.t3510 VSS.t2040 1551.14
R6994 VSS.t1238 VSS.t4328 1551.14
R6995 VSS.t3895 VSS.t3355 1551.14
R6996 VSS.t2391 VSS.t1246 1551.14
R6997 VSS.t4340 VSS.t3872 1551.14
R6998 VSS.t2524 VSS.t3525 1551.14
R6999 VSS.t1342 VSS.t2057 1551.14
R7000 VSS.t2227 VSS.t1183 1551.14
R7001 VSS.t2059 VSS.t2227 1551.14
R7002 VSS.t1185 VSS.t2379 1551.14
R7003 VSS.t2293 VSS.t1707 1551.14
R7004 VSS.t3206 VSS.t1653 1551.14
R7005 VSS.t3444 VSS.t2110 1551.14
R7006 VSS.t3249 VSS.t2276 1551.14
R7007 VSS.t1495 VSS.t3149 1551.14
R7008 VSS.t1873 VSS.t1293 1551.14
R7009 VSS.t3267 VSS.t2032 1551.14
R7010 VSS.t3267 VSS.t1289 1551.14
R7011 VSS.t3906 VSS.t2167 1551.14
R7012 VSS.t3245 VSS.t3563 1551.14
R7013 VSS.t1300 VSS.t1505 1551.14
R7014 VSS.t3860 VSS.t3953 1551.14
R7015 VSS.t4124 VSS.t3408 1551.14
R7016 VSS.t928 VSS.t2886 1551.14
R7017 VSS.t3854 VSS.t1757 1551.14
R7018 VSS.t2504 VSS.t4277 1551.14
R7019 VSS.t4277 VSS.t2548 1551.14
R7020 VSS.t1460 VSS.t1419 1551.14
R7021 VSS.t3402 VSS.t3426 1551.14
R7022 VSS.t2246 VSS.t3231 1551.14
R7023 VSS.t1236 VSS.t1232 1551.14
R7024 VSS.t2139 VSS.t2552 1551.14
R7025 VSS.t1464 VSS.t3255 1551.14
R7026 VSS.t2491 VSS.t3087 1551.14
R7027 VSS.t2584 VSS.t3972 1551.14
R7028 VSS.t4128 VSS.t2584 1551.14
R7029 VSS.t1992 VSS.t1533 1551.14
R7030 VSS.t1029 VSS.t2999 1551.14
R7031 VSS.t3566 VSS.t3210 1551.14
R7032 VSS.t3229 VSS.t3752 1551.14
R7033 VSS.t3166 VSS.t965 1551.14
R7034 VSS.t3122 VSS.t2535 1551.14
R7035 VSS.t1392 VSS.t973 1551.14
R7036 VSS.t4095 VSS.t2180 1551.14
R7037 VSS.t3886 VSS.t1529 1551.14
R7038 VSS.t3726 VSS.t3694 1551.14
R7039 VSS.t4231 VSS.t2898 1551.14
R7040 VSS.t1261 VSS.t1212 1551.14
R7041 VSS.t1278 VSS.t3100 1551.14
R7042 VSS.t3189 VSS.t3949 1551.14
R7043 VSS.t2334 VSS.t4321 1551.14
R7044 VSS.t2906 VSS.t2334 1551.14
R7045 VSS.t3032 VSS.t4251 1551.14
R7046 VSS.t985 VSS.t1139 1551.14
R7047 VSS.t1638 VSS.t1473 1551.14
R7048 VSS.t2957 VSS.t954 1551.14
R7049 VSS.t1987 VSS.t2468 1551.14
R7050 VSS.t2322 VSS.t1000 1551.14
R7051 VSS.t1387 VSS.t1291 1551.14
R7052 VSS.t1550 VSS.t2233 1551.14
R7053 VSS.t1295 VSS.t1550 1551.14
R7054 VSS.t2286 VSS.t2493 1551.14
R7055 VSS.t1983 VSS.t2900 1551.14
R7056 VSS.t2827 VSS.t3038 1551.14
R7057 VSS.t3457 VSS.t4216 1551.14
R7058 VSS.t2770 VSS.t1634 1551.14
R7059 VSS.t2657 VSS.t3451 1551.14
R7060 VSS.t1586 VSS.t2159 1551.14
R7061 VSS.t4044 VSS.t4018 1551.14
R7062 VSS.t2965 VSS.t4044 1551.14
R7063 VSS.t3935 VSS.t2604 1551.14
R7064 VSS.t2016 VSS.t2973 1551.14
R7065 VSS.t1715 VSS.t3924 1551.14
R7066 VSS.t3251 VSS.t956 1551.14
R7067 VSS.t3285 VSS.t3488 1551.14
R7068 VSS.t3931 VSS.t2607 1551.14
R7069 VSS.t1151 VSS.t2694 1551.14
R7070 VSS.t4024 VSS.t2835 1551.14
R7071 VSS.t2284 VSS.t1477 1551.14
R7072 VSS.t2554 VSS.t3891 1551.14
R7073 VSS.t2163 VSS.t2952 1551.14
R7074 VSS.t2961 VSS.t3625 1551.14
R7075 VSS.t2466 VSS.t3464 1551.14
R7076 VSS.t2346 VSS.t3762 1551.14
R7077 VSS.t2633 VSS.t1177 1551.14
R7078 VSS.t2288 VSS.t3550 1551.14
R7079 VSS.t1755 VSS.t2526 1551.14
R7080 VSS.t3389 VSS.t2182 1551.14
R7081 VSS.t1143 VSS.t3627 1551.14
R7082 VSS.t4151 VSS.t2211 1551.14
R7083 VSS.t2772 VSS.t3118 1551.14
R7084 VSS.t3959 VSS.t4275 1551.14
R7085 VSS.t3959 VSS.t3334 1551.14
R7086 VSS.t3963 VSS.t1852 1551.14
R7087 VSS.t1918 VSS.t1336 1551.14
R7088 VSS.t4176 VSS.t3018 1551.14
R7089 VSS.t2063 VSS.t1251 1551.14
R7090 VSS.t1770 VSS.t3338 1551.14
R7091 VSS.t1405 VSS.t2131 1551.14
R7092 VSS.t3083 VSS.t1226 1551.14
R7093 VSS.t3712 VSS.t4336 1551.14
R7094 VSS.t4336 VSS.t3233 1551.14
R7095 VSS.t2711 VSS.t2069 1551.14
R7096 VSS.t2042 VSS.t2118 1551.14
R7097 VSS.t1763 VSS.t4241 1551.14
R7098 VSS.t3073 VSS.t1021 1551.14
R7099 VSS.t2963 VSS.t3561 1551.14
R7100 VSS.t1807 VSS.t4355 1551.14
R7101 VSS.t2785 VSS.t1374 1551.14
R7102 VSS.t2938 VSS.t3728 1551.14
R7103 VSS.t3728 VSS.t2594 1551.14
R7104 VSS.t1033 VSS.t3241 1551.14
R7105 VSS.t4122 VSS.t3484 1551.14
R7106 VSS.t2462 VSS.t1458 1551.14
R7107 VSS.t1940 VSS.t3519 1551.14
R7108 VSS.t1914 VSS.t3440 1551.14
R7109 VSS.t1772 VSS.t3181 1551.14
R7110 VSS.t2478 VSS.t2328 1551.14
R7111 VSS.t4077 VSS.t1242 1551.14
R7112 VSS.t2307 VSS.t1306 1551.14
R7113 VSS.t3554 VSS.t2894 1551.14
R7114 VSS.t2235 VSS.t2720 1551.14
R7115 VSS.t2448 VSS.t4350 1551.14
R7116 VSS.t1214 VSS.t2971 1551.14
R7117 VSS.t3047 VSS.t3067 1551.14
R7118 VSS.t3191 VSS.t2870 1551.14
R7119 VSS.t2402 VSS.t2724 1551.14
R7120 VSS.t3324 VSS.t2402 1551.14
R7121 VSS.t2146 VSS.t4239 1551.14
R7122 VSS.t1774 VSS.t952 1551.14
R7123 VSS.t3916 VSS.t3521 1551.14
R7124 VSS.t3417 VSS.t3649 1551.14
R7125 VSS.t3411 VSS.t2702 1551.14
R7126 VSS.t1881 VSS.t1002 1551.14
R7127 VSS.t2969 VSS.t1297 1551.14
R7128 VSS.t2829 VSS.t2258 1551.14
R7129 VSS.t1421 VSS.t2829 1551.14
R7130 VSS.t1253 VSS.t2934 1551.14
R7131 VSS.t3714 VSS.t4297 1551.14
R7132 VSS.t3615 VSS.t3740 1551.14
R7133 VSS.t3462 VSS.t3793 1551.14
R7134 VSS.t3672 VSS.t3077 1551.14
R7135 VSS.t2696 VSS.t2540 1551.14
R7136 VSS.t2508 VSS.t3094 1551.14
R7137 VSS.t2120 VSS.t1244 1551.14
R7138 VSS.t2831 VSS.n972 1551.14
R7139 VSS.t4283 VSS.t1590 1551.14
R7140 VSS.t3508 VSS.t1515 1551.14
R7141 VSS.t2866 VSS.t4005 1551.14
R7142 VSS.t1614 VSS.t1031 1551.14
R7143 VSS.t960 VSS.t2622 1551.14
R7144 VSS.t4287 VSS.t3750 1551.14
R7145 VSS.t3843 VSS.t1651 1551.14
R7146 VSS.t3843 VSS.t2202 1551.14
R7147 VSS.t1705 VSS.t3664 1551.14
R7148 VSS.t3043 VSS.t2200 1551.14
R7149 VSS.t2510 VSS.t3623 1551.14
R7150 VSS.t1481 VSS.t1548 1551.14
R7151 VSS.t1608 VSS.t3533 1551.14
R7152 VSS.t3644 VSS.t3841 1551.14
R7153 VSS.t3243 VSS.t2631 1551.14
R7154 VSS.t2165 VSS.t967 1551.14
R7155 VSS.t4051 VSS.t2282 1551.14
R7156 VSS.t2546 VSS.t979 1551.14
R7157 VSS.t3834 VSS.t1964 1551.14
R7158 VSS.t2018 VSS.t3177 1551.14
R7159 VSS.t3552 VSS.t2157 1551.14
R7160 VSS.t1588 VSS.t3145 1551.14
R7161 VSS.t4120 VSS.t1027 1551.14
R7162 VSS.t1759 VSS.t3678 1551.14
R7163 VSS.t2803 VSS.t1179 1551.14
R7164 VSS.t3506 VSS.t3153 1551.14
R7165 VSS.t3272 VSS.t3619 1551.14
R7166 VSS.t2728 VSS.t4243 1551.14
R7167 VSS.t1200 VSS.t3582 1551.14
R7168 VSS.t3253 VSS.t3024 1551.14
R7169 VSS.t3253 VSS.t4022 1551.14
R7170 VSS.t3014 VSS.t3393 1551.14
R7171 VSS.t2698 VSS.t2908 1551.14
R7172 VSS.t2730 VSS.t1662 1551.14
R7173 VSS.t4028 VSS.t4069 1551.14
R7174 VSS.t4016 VSS.t3884 1551.14
R7175 VSS.t4172 VSS.t3710 1551.14
R7176 VSS.t2569 VSS.t3326 1551.14
R7177 VSS.t3764 VSS.t2955 1551.14
R7178 VSS.t2955 VSS.t2350 1551.14
R7179 VSS.t3850 VSS.t2833 1551.14
R7180 VSS.t4301 VSS.t3459 1551.14
R7181 VSS.t2783 VSS.t2936 1551.14
R7182 VSS.t2389 VSS.t2359 1551.14
R7183 VSS.t3235 VSS.t2777 1551.14
R7184 VSS.t2148 VSS.t4093 1551.14
R7185 VSS.t2851 VSS.t4010 1551.14
R7186 VSS.t2902 VSS.t3287 1551.14
R7187 VSS.t3287 VSS.t2102 1551.14
R7188 VSS.t975 VSS.t3453 1551.14
R7189 VSS.t191 VSS.t234 1551.14
R7190 VSS.t3937 VSS.t3817 1551.14
R7191 VSS.t1396 VSS.t2882 1551.14
R7192 VSS.t4344 VSS.t2932 1551.14
R7193 VSS.t1544 VSS.t1145 1551.14
R7194 VSS.t3227 VSS.t1648 1551.14
R7195 VSS.t2857 VSS.t3353 1551.14
R7196 VSS.t2444 VSS.t3223 1551.14
R7197 VSS.t3160 VSS.t2444 1551.14
R7198 VSS.t1713 VSS.t3617 1551.14
R7199 VSS.t2330 VSS.t2736 1551.14
R7200 VSS.t2332 VSS.t3237 1551.14
R7201 VSS.t1539 VSS.t1916 1551.14
R7202 VSS.t3302 VSS.t3089 1551.14
R7203 VSS.t1281 VSS.t1467 1551.14
R7204 VSS.t3363 VSS.t2718 1551.14
R7205 VSS.t1423 VSS.t3826 1551.14
R7206 VSS.t2204 VSS.t1423 1551.14
R7207 VSS.t2615 VSS.t1885 1551.14
R7208 VSS.t3722 VSS.t3660 1551.14
R7209 VSS.t3349 VSS.t3922 1551.14
R7210 VSS.t3965 VSS.t2175 1551.14
R7211 VSS.t4271 VSS.t3102 1551.14
R7212 VSS.t3468 VSS.t4067 1551.14
R7213 VSS.t2876 VSS.t3304 1551.14
R7214 VSS.t2355 VSS.t1893 1551.14
R7215 VSS.t2381 VSS.t3832 1551.14
R7216 VSS.t4332 VSS.t2197 1551.14
R7217 VSS.t3423 VSS.t2100 1551.14
R7218 VSS.t3142 VSS.t4279 1551.14
R7219 VSS.t3535 VSS.t3413 1551.14
R7220 VSS.t1469 VSS.t1338 1551.14
R7221 VSS.t1019 VSS.t3662 1551.14
R7222 VSS.t1019 VSS.t2418 1551.14
R7223 VSS.t1499 VSS.t3085 1551.14
R7224 VSS.t1930 VSS.t4257 1551.14
R7225 VSS.t3264 VSS.t3185 1551.14
R7226 VSS.t2446 VSS.t1326 1551.14
R7227 VSS.t4178 VSS.t2456 1551.14
R7228 VSS.t3601 VSS.t3225 1551.14
R7229 VSS.t1920 VSS.t4145 1551.14
R7230 VSS.t3893 VSS.t1425 1551.14
R7231 VSS.t2625 VSS.t2726 1551.14
R7232 VSS.t3880 VSS.t2896 1551.14
R7233 VSS.t1409 VSS.t2940 1551.14
R7234 VSS.t1616 VSS.t4149 1551.14
R7235 VSS.t1666 VSS.t1136 1551.14
R7236 VSS.t2644 VSS.t2704 1551.14
R7237 VSS.t3391 VSS.t1283 1551.14
R7238 VSS.t2892 VSS.t2239 1551.14
R7239 VSS.t4338 VSS.t2984 1551.14
R7240 VSS.t1134 VSS.t2104 1551.14
R7241 VSS.t2085 VSS.t1394 1551.14
R7242 VSS.t2528 VSS.t1497 1551.14
R7243 VSS.t2486 VSS.t4020 1551.14
R7244 VSS.t3080 VSS.t2000 1551.14
R7245 VSS.t3080 VSS.t2967 1551.14
R7246 VSS.t3173 VSS.t3274 1551.14
R7247 VSS.t3967 VSS.t2071 1551.14
R7248 VSS.t4227 VSS.t3939 1551.14
R7249 VSS.t3217 VSS.t2408 1551.14
R7250 VSS.t2506 VSS.t3016 1551.14
R7251 VSS.t1189 VSS.t3478 1551.14
R7252 VSS.t2618 VSS.t3807 1551.14
R7253 VSS.t2116 VSS.t4255 1551.14
R7254 VSS.t2847 VSS.t4237 1551.14
R7255 VSS.t2264 VSS.t4233 1551.14
R7256 VSS.t2357 VSS.t3208 1551.14
R7257 VSS.t1584 VSS.t2133 1551.14
R7258 VSS.t1610 VSS.t3870 1551.14
R7259 VSS.t2482 VSS.t1259 1551.14
R7260 VSS.t2209 VSS.t1443 1551.14
R7261 VSS.t2819 VSS.t4330 1551.14
R7262 VSS.t2067 VSS.t1658 1551.14
R7263 VSS.t3782 VSS.t3336 1551.14
R7264 VSS.t2191 VSS.t3215 1551.14
R7265 VSS.t2250 VSS.n1329 1551.14
R7266 VSS.t4026 VSS.t2563 1551.14
R7267 VSS.t3257 VSS.t2225 1551.14
R7268 VSS.t3120 VSS.t3819 1551.14
R7269 VSS.t3912 VSS.t3612 1551.14
R7270 VSS.t3547 VSS.t2458 1551.14
R7271 VSS.t1664 VSS.t3647 1551.14
R7272 VSS.t2740 VSS.t3997 1551.14
R7273 VSS.t3179 VSS.t3920 1551.14
R7274 VSS.t3179 VSS.t2565 1551.14
R7275 VSS.t3395 VSS.t1564 1551.14
R7276 VSS.t3951 VSS.t3957 1551.14
R7277 VSS.t1194 VSS.t3995 1551.14
R7278 VSS.t1962 VSS.t2734 1551.14
R7279 VSS.t3605 VSS.t2141 1551.14
R7280 VSS.t1224 VSS.t1612 1551.14
R7281 VSS.t3164 VSS.t1162 1551.14
R7282 VSS.t4065 VSS.t2653 1551.14
R7283 VSS.t1240 VSS.t2978 1551.14
R7284 VSS.t4071 VSS.t4130 1551.14
R7285 VSS.t2868 VSS.t2237 1551.14
R7286 VSS.t335 VSS.t1314 1551.14
R7287 VSS.t770 VSS.t820 1551.14
R7288 VSS.t3480 VSS.t1181 1551.14
R7289 VSS.t1632 VSS.t2412 1551.14
R7290 VSS.t4055 VSS.t4324 1551.14
R7291 VSS.t971 VSS.t3610 1551.14
R7292 VSS.t3852 VSS.t2460 1551.14
R7293 VSS.t4346 VSS.t2112 1551.14
R7294 VSS.n1451 VSS.t2533 1551.14
R7295 VSS.t2815 VSS.t15 1551.14
R7296 VSS.t816 VSS.t1868 1551.14
R7297 VSS.n1430 VSS.t3293 1551.14
R7298 VSS.t3383 VSS.t4210 1551.14
R7299 VSS.n927 VSS.t1912 1528.05
R7300 VSS.t1257 VSS.t2244 1523.44
R7301 VSS.t1700 VSS.t4299 1523.44
R7302 VSS.n1994 VSS.t1075 1514.2
R7303 VSS.t1017 VSS.t4303 1495.74
R7304 VSS.t1379 VSS.t2173 1495.74
R7305 VSS.t11 VSS.t2744 1486.51
R7306 VSS.t1578 VSS.t1875 1481.89
R7307 VSS.t4112 VSS.t1946 1481.89
R7308 VSS.t4034 VSS.t287 1444.96
R7309 VSS.n2537 VSS.n2536 1443.52
R7310 VSS.t4073 VSS.t2152 1440.34
R7311 VSS.t141 VSS.t1255 1440.34
R7312 VSS.t489 VSS.t1535 1440.34
R7313 VSS.t1554 VSS.t4115 1440.34
R7314 VSS.t1487 VSS.t3595 1440.34
R7315 VSS.t1867 VSS.t2821 1440.34
R7316 VSS.t4036 VSS.t4003 1440.34
R7317 VSS.t2982 VSS.t1485 1440.34
R7318 VSS.n436 VSS.t3734 1435.72
R7319 VSS.n2432 VSS.n2431 1432.24
R7320 VSS.t3736 VSS.t3442 1426.49
R7321 VSS.t833 VSS.t2416 1412.64
R7322 VSS.t678 VSS.t114 1403.41
R7323 VSS.t3214 VSS.t1815 1398.79
R7324 VSS.t2243 VSS.t2864 1398.79
R7325 VSS.t4220 VSS.t2008 1398.79
R7326 VSS.n399 VSS.t845 1398.79
R7327 VSS.t2880 VSS.t3110 1389.56
R7328 VSS.n2538 VSS.n2537 1387.96
R7329 VSS.t514 VSS.t2336 1384.94
R7330 VSS.t2682 VSS.n72 1384.94
R7331 VSS.t2684 VSS.n70 1384.94
R7332 VSS.t2676 VSS.n69 1384.94
R7333 VSS.t682 VSS.n68 1384.94
R7334 VSS.t404 VSS.n67 1384.94
R7335 VSS.t394 VSS.n66 1384.94
R7336 VSS.n575 VSS.t402 1384.94
R7337 VSS.t685 VSS.t1489 1366.48
R7338 VSS.t4187 VSS.t4334 1366.48
R7339 VSS.t4139 VSS.t4008 1366.48
R7340 VSS.t4197 VSS.t996 1366.48
R7341 VSS.t990 VSS.t327 1366.48
R7342 VSS.t2005 VSS.t525 1366.48
R7343 VSS.t2484 VSS.t4186 1366.48
R7344 VSS.t1210 VSS.t1895 1366.48
R7345 VSS.t352 VSS.n636 1366.48
R7346 VSS.n419 VSS.t408 1366.48
R7347 VSS.n552 VSS.t846 1366.48
R7348 VSS.t3187 VSS.t924 1366.48
R7349 VSS.t4089 VSS.t3779 1361.86
R7350 VSS.n2422 VSS.t208 1335.3
R7351 VSS.t3361 VSS.t2888 1334.16
R7352 VSS.t915 VSS.n459 1332.99
R7353 VSS.t1111 VSS.t645 1329.55
R7354 VSS.n2219 VSS.n2218 1322.26
R7355 VSS.n2220 VSS.n2219 1322.26
R7356 VSS.n2221 VSS.n2220 1322.26
R7357 VSS.n2222 VSS.n2221 1322.26
R7358 VSS.n2223 VSS.n2222 1322.26
R7359 VSS.n2224 VSS.n2223 1322.26
R7360 VSS.n2225 VSS.n2224 1322.26
R7361 VSS.n2226 VSS.n2225 1322.26
R7362 VSS.n2227 VSS.n2226 1322.26
R7363 VSS.n2228 VSS.n2227 1322.26
R7364 VSS.n2229 VSS.n2228 1322.26
R7365 VSS.n2230 VSS.n2229 1322.26
R7366 VSS.n2231 VSS.n2230 1322.26
R7367 VSS.n459 VSS.t396 1319.62
R7368 VSS.n764 VSS.t4320 1311.08
R7369 VSS.t2924 VSS.t3063 1297.23
R7370 VSS.t2279 VSS.t2746 1297.23
R7371 VSS.t2171 VSS.t2470 1288
R7372 VSS.n984 VSS.t1514 1274.15
R7373 VSS.n644 VSS.t2879 1274.15
R7374 VSS.t3401 VSS.t3738 1269.53
R7375 VSS.t189 VSS.t1956 1260.3
R7376 VSS.n2433 VSS.n2432 1242.47
R7377 VSS.t3322 VSS.t2122 1241.83
R7378 VSS.n2440 VSS.n2439 1238.48
R7379 VSS.t831 VSS.t4269 1237.22
R7380 VSS.t1377 VSS.t1765 1237.22
R7381 VSS.t3406 VSS.t1813 1237.22
R7382 VSS.t4223 VSS.t2558 1237.22
R7383 VSS.t4059 VSS.t2038 1237.22
R7384 VSS.t540 VSS.t478 1237.22
R7385 VSS.t899 VSS.t1304 1237.22
R7386 VSS.t1207 VSS.t2801 1237.22
R7387 VSS.t1068 VSS.t1285 1237.22
R7388 VSS.t708 VSS.t1081 1236.7
R7389 VSS.t3955 VSS.t1902 1227.98
R7390 VSS.t3688 VSS.t1856 1227.98
R7391 VSS.t2489 VSS.t544 1218.75
R7392 VSS.t2073 VSS.n774 1218.75
R7393 VSS.t10 VSS.n1458 1218.75
R7394 VSS.t3556 VSS.t128 1214.13
R7395 VSS.t1306 VSS.t3789 1200.28
R7396 VSS.t2579 VSS.t523 1200.28
R7397 VSS.t1519 VSS.t3587 1200.28
R7398 VSS.t2038 VSS.t4285 1200.28
R7399 VSS.t1767 VSS.t494 1200.28
R7400 VSS.t1274 VSS.t3381 1200.28
R7401 VSS.t806 VSS.t1802 1200.28
R7402 VSS.t2496 VSS.t3158 1200.28
R7403 VSS.t1023 VSS.t804 1200.28
R7404 VSS.t1299 VSS.t819 1186.43
R7405 VSS.t523 VSS.t1711 1181.82
R7406 VSS.t521 VSS.t2127 1181.82
R7407 VSS.t482 VSS.t1646 1181.82
R7408 VSS.t789 VSS.t1580 1181.82
R7409 VSS.t505 VSS.t1035 1181.82
R7410 VSS.t4247 VSS.t810 1181.82
R7411 VSS.t1198 VSS.t783 1181.82
R7412 VSS.t2296 VSS.t325 1181.82
R7413 VSS.t763 VSS.t3428 1181.82
R7414 VSS.t793 VSS.t3732 1181.82
R7415 VSS.t827 VSS.t3690 1181.82
R7416 VSS.t3112 VSS.t2586 1181.82
R7417 VSS.t835 VSS.t1070 1181.82
R7418 VSS.t1087 VSS.t4253 1172.59
R7419 VSS.t1249 VSS.t3927 1167.97
R7420 VSS.t2003 VSS.t1954 1167.97
R7421 VSS.t494 VSS.t1216 1167.97
R7422 VSS.t535 VSS.t2994 1167.97
R7423 VSS.t542 VSS.t3746 1167.97
R7424 VSS.n1995 VSS.t3279 1149.5
R7425 VSS.t1417 VSS.t3010 1149.5
R7426 VSS.t1989 VSS.t4059 1144.89
R7427 VSS.t4191 VSS.t1501 1140.27
R7428 VSS.t3708 VSS.t3196 1131.04
R7429 VSS.t4206 VSS.t2775 1126.42
R7430 VSS.t2879 VSS.t285 1126.42
R7431 VSS.t1158 VSS.t4012 1126.42
R7432 VSS.t3529 VSS.t3471 1121.8
R7433 VSS.n788 VSS.t1166 1112.57
R7434 VSS.t2843 VSS.t4221 1112.57
R7435 VSS.t3202 VSS.t1507 1103.34
R7436 VSS.t935 VSS.t3760 1103.34
R7437 VSS.t684 VSS.t4038 1103.34
R7438 VSS.n655 VSS.t2320 1103.34
R7439 VSS.t3874 VSS.t694 1089.49
R7440 VSS.t1906 VSS.t3668 1089.49
R7441 VSS.t4320 VSS.t289 1089.49
R7442 VSS.t4091 VSS.t7 1089.49
R7443 VSS.t3061 VSS.t513 1089.49
R7444 VSS.t3320 VSS.t3874 1084.87
R7445 VSS.t4147 VSS.t1132 1084.87
R7446 VSS.t2229 VSS.t1039 1080.26
R7447 VSS.t2476 VSS.t2090 1071.02
R7448 VSS.t1650 VSS.t2254 1071.02
R7449 VSS.t2862 VSS.t3948 1071.02
R7450 VSS.n1852 VSS.t2998 1066.41
R7451 VSS.t958 VSS.t681 1066.41
R7452 VSS.t837 VSS.t3075 1066.41
R7453 VSS.t3283 VSS.t1650 1066.41
R7454 VSS.t2538 VSS.t2156 1061.79
R7455 VSS.n1717 VSS.t2655 1052.56
R7456 VSS.t779 VSS.n856 1052.56
R7457 VSS.n2425 VSS.n2424 1048.71
R7458 VSS.t1980 VSS.t2050 1047.94
R7459 VSS.t44 VSS.t542 1047.94
R7460 VSS.t796 VSS.t2268 1047.67
R7461 VSS.t2035 VSS.t2742 1038.71
R7462 VSS.t2108 VSS.t2890 1038.71
R7463 VSS.t4087 VSS.t3560 1038.71
R7464 VSS.t3766 VSS.t2275 1038.71
R7465 VSS.t3030 VSS.t3579 1038.71
R7466 VSS.t1592 VSS.t3642 1038.71
R7467 VSS.t3066 VSS.t1900 1038.71
R7468 VSS.t2817 VSS.t3096 1038.71
R7469 VSS.t3690 VSS.t2588 1038.71
R7470 VSS.t1562 VSS.t3947 1038.71
R7471 VSS.n1023 VSS.t992 1034.09
R7472 VSS.t1089 VSS.n1023 1034.09
R7473 VSS.t1668 VSS.t947 1034.09
R7474 VSS.t947 VSS.t1692 1034.09
R7475 VSS.t4305 VSS.t4311 1034.09
R7476 VSS.t4309 VSS.t4307 1034.09
R7477 VSS.t1042 VSS.t1056 1034.09
R7478 VSS.t1050 VSS.t1048 1034.09
R7479 VSS.t1054 VSS.t1044 1034.09
R7480 VSS.t1046 VSS.t1052 1034.09
R7481 VSS.t1729 VSS.t1721 1034.09
R7482 VSS.t1717 VSS.t1727 1034.09
R7483 VSS.t1725 VSS.t1731 1034.09
R7484 VSS.t1723 VSS.t1719 1034.09
R7485 VSS.t787 VSS.t771 1034.09
R7486 VSS.t771 VSS.t695 1034.09
R7487 VSS.t3590 VSS.t2515 1034.09
R7488 VSS.t2375 VSS.t2367 1034.09
R7489 VSS.t2373 VSS.t2363 1034.09
R7490 VSS.t2377 VSS.t2369 1034.09
R7491 VSS.t2808 VSS.t529 1034.09
R7492 VSS.t2810 VSS.t2808 1034.09
R7493 VSS.t2680 VSS.t2036 1034.09
R7494 VSS.t3813 VSS.t1850 1034.09
R7495 VSS.t1598 VSS.t1952 1034.09
R7496 VSS.t1952 VSS.t1602 1034.09
R7497 VSS.t1602 VSS.t2079 1034.09
R7498 VSS.t1990 VSS.t1600 1034.09
R7499 VSS.n912 VSS.t3311 1034.09
R7500 VSS.t3538 VSS.n912 1034.09
R7501 VSS.t2410 VSS.t3538 1034.09
R7502 VSS.t1456 VSS.t2410 1034.09
R7503 VSS.t2348 VSS.t1456 1034.09
R7504 VSS.t1863 VSS.t2348 1034.09
R7505 VSS.t2797 VSS.t1863 1034.09
R7506 VSS.t1537 VSS.t2797 1034.09
R7507 VSS.t3344 VSS.t1537 1034.09
R7508 VSS.t2853 VSS.t3344 1034.09
R7509 VSS.t2706 VSS.t2853 1034.09
R7510 VSS.t2385 VSS.t2706 1034.09
R7511 VSS.t1813 VSS.t283 1034.09
R7512 VSS.t1811 VSS.t1471 1034.09
R7513 VSS.t1568 VSS.t1761 1034.09
R7514 VSS.t2216 VSS.t1606 1034.09
R7515 VSS.t4281 VSS.t3575 1034.09
R7516 VSS.t2910 VSS.t1561 1034.09
R7517 VSS.t2922 VSS.t3270 1034.09
R7518 VSS.t3797 VSS.t959 1034.09
R7519 VSS.t508 VSS.t191 1034.09
R7520 VSS.t1747 VSS.t1753 1034.09
R7521 VSS.t307 VSS.t313 1034.09
R7522 VSS.t4133 VSS.t420 1034.09
R7523 VSS.t470 VSS.t423 1034.09
R7524 VSS.n871 VSS.t2229 1034.09
R7525 VSS.t1955 VSS.t3449 1034.09
R7526 VSS.t3449 VSS.t2262 1034.09
R7527 VSS.t1138 VSS.t3571 1034.09
R7528 VSS.n781 VSS.t4143 1034.09
R7529 VSS.t1479 VSS.n781 1034.09
R7530 VSS.t863 VSS.t867 1034.09
R7531 VSS.t301 VSS.t297 1034.09
R7532 VSS.t291 VSS.t301 1034.09
R7533 VSS.t295 VSS.t291 1034.09
R7534 VSS.t303 VSS.t305 1034.09
R7535 VSS.t3945 VSS.t3946 1034.09
R7536 VSS.t2601 VSS.t3171 1034.09
R7537 VSS.t3584 VSS.t422 1034.09
R7538 VSS.t2361 VSS.t507 1034.09
R7539 VSS.t48 VSS.t426 1034.09
R7540 VSS.t46 VSS.t50 1034.09
R7541 VSS.t1897 VSS.t1012 1034.09
R7542 VSS.t2077 VSS.t2075 1034.09
R7543 VSS.t159 VSS.t161 1034.09
R7544 VSS.t147 VSS.t145 1034.09
R7545 VSS.t149 VSS.t143 1034.09
R7546 VSS.t169 VSS.t153 1034.09
R7547 VSS.t2047 VSS.t1888 1034.09
R7548 VSS.t3140 VSS.t1340 1034.09
R7549 VSS.t711 VSS.t702 1034.09
R7550 VSS.t2668 VSS.t2690 1034.09
R7551 VSS.t2662 VSS.t2664 1034.09
R7552 VSS.t1553 VSS.t969 1034.09
R7553 VSS.t1555 VSS.t2672 1034.09
R7554 VSS.t2672 VSS.t1103 1034.09
R7555 VSS.t1103 VSS.t682 1034.09
R7556 VSS.t398 VSS.t358 1034.09
R7557 VSS.t333 VSS.t364 1034.09
R7558 VSS.t1376 VSS.t3585 1034.09
R7559 VSS.t3580 VSS.t404 1034.09
R7560 VSS.t4046 VSS.t1566 1034.09
R7561 VSS.t1985 VSS.t4046 1034.09
R7562 VSS.t3651 VSS.t1985 1034.09
R7563 VSS.t2781 VSS.t3651 1034.09
R7564 VSS.t3638 VSS.t2781 1034.09
R7565 VSS.t3929 VSS.t3638 1034.09
R7566 VSS.t3332 VSS.t3929 1034.09
R7567 VSS.t2326 VSS.t3332 1034.09
R7568 VSS.t2098 VSS.t2326 1034.09
R7569 VSS.t1493 VSS.t2098 1034.09
R7570 VSS.t2700 VSS.t1493 1034.09
R7571 VSS.t3247 VSS.t2700 1034.09
R7572 VSS.t1703 VSS.t3247 1034.09
R7573 VSS.t3262 VSS.t1703 1034.09
R7574 VSS.t2986 VSS.t3262 1034.09
R7575 VSS.t4164 VSS.t4168 1034.09
R7576 VSS.t4160 VSS.t4166 1034.09
R7577 VSS.t4156 VSS.t4170 1034.09
R7578 VSS.t879 VSS.t877 1034.09
R7579 VSS.t883 VSS.t871 1034.09
R7580 VSS.t885 VSS.t873 1034.09
R7581 VSS.t650 VSS.t658 1034.09
R7582 VSS.t23 VSS.t131 1034.09
R7583 VSS.t2320 VSS.t1390 1034.09
R7584 VSS.t609 VSS.t611 1034.09
R7585 VSS.t905 VSS.t913 1034.09
R7586 VSS.t649 VSS.t652 1034.09
R7587 VSS.t1315 VSS.t3069 1034.09
R7588 VSS.t2014 VSS.t3371 1034.09
R7589 VSS.t2303 VSS.t2732 1034.09
R7590 VSS.t3065 VSS.t3385 1034.09
R7591 VSS.t2298 VSS.t4323 1034.09
R7592 VSS.t3346 VSS.t1503 1034.09
R7593 VSS.t4104 VSS.t2818 1034.09
R7594 VSS.t1488 VSS.t1527 1034.09
R7595 VSS.t1684 VSS.t1678 1034.09
R7596 VSS.t1682 VSS.t1670 1034.09
R7597 VSS.t661 VSS.t643 1034.09
R7598 VSS.t4 VSS.t663 1034.09
R7599 VSS.t472 VSS.t4 1034.09
R7600 VSS.t464 VSS.t472 1034.09
R7601 VSS.t555 VSS.t464 1034.09
R7602 VSS.t36 VSS.t32 1034.09
R7603 VSS.t42 VSS.t40 1034.09
R7604 VSS.t922 VSS.t926 1034.09
R7605 VSS.t920 VSS.t922 1034.09
R7606 VSS.n1516 VSS.t2639 1034.09
R7607 VSS.t1870 VSS.t3961 1034.09
R7608 VSS.t175 VSS.t173 1034.09
R7609 VSS.t4263 VSS.t4265 1034.09
R7610 VSS.t4037 VSS.t1640 1034.09
R7611 VSS.t2586 VSS.t406 1034.09
R7612 VSS.t3770 VSS.t3772 1034.09
R7613 VSS.t328 VSS.t753 1034.09
R7614 VSS.t4042 VSS.t1415 1034.09
R7615 VSS.t3876 VSS.t2344 1034.09
R7616 VSS.t2301 VSS.t2477 1034.09
R7617 VSS.t2012 VSS.t2299 1034.09
R7618 VSS.t981 VSS.n631 1034.09
R7619 VSS.n631 VSS.t2799 1034.09
R7620 VSS.t3706 VSS.t3704 1034.09
R7621 VSS.t2027 VSS.t655 1034.09
R7622 VSS.t3470 VSS.t3109 1034.09
R7623 VSS.t930 VSS.t466 1034.09
R7624 VSS.t2975 VSS.t1562 1034.09
R7625 VSS.t1109 VSS.t19 1034.09
R7626 VSS.t3342 VSS.t3340 1034.09
R7627 VSS.t847 VSS.t370 1034.09
R7628 VSS.t1128 VSS.t847 1034.09
R7629 VSS.t2452 VSS.t3404 1034.09
R7630 VSS.t1310 VSS.t551 1029.47
R7631 VSS.t2207 VSS.t2295 1029.47
R7632 VSS.t1058 VSS.t1218 1020.24
R7633 VSS.t1879 VSS.t1627 1020.24
R7634 VSS.t496 VSS.t1101 1020.24
R7635 VSS.t1936 VSS.t2992 1020.24
R7636 VSS.t3633 VSS.t3748 1020.24
R7637 VSS.t3369 VSS.t187 1020.24
R7638 VSS.t4074 VSS.n915 1015.62
R7639 VSS.t2155 VSS.n921 1015.62
R7640 VSS.t4031 VSS.t1220 1015.62
R7641 VSS.n774 VSS.t163 1015.62
R7642 VSS.t3824 VSS.t4164 1015.62
R7643 VSS.t1806 VSS.t2990 1015.62
R7644 VSS.t3435 VSS.t3742 1015.62
R7645 VSS.t2550 VSS.n390 1015.62
R7646 VSS.t1011 VSS.t183 1015.62
R7647 VSS.t2799 VSS.t1743 1015.62
R7648 VSS.t2512 VSS.t2624 1011.01
R7649 VSS.n2549 VSS.n11 1007.82
R7650 VSS.t4140 VSS.t3156 1006.39
R7651 VSS.t3658 VSS.t2613 1006.39
R7652 VSS.t3004 VSS.t3002 1006.39
R7653 VSS.t3882 VSS.t1318 1006.39
R7654 VSS.t3151 VSS.t2314 1001.78
R7655 VSS.t1944 VSS.t4289 997.159
R7656 VSS.t3026 VSS.t232 997.159
R7657 VSS.t4348 VSS.t1263 997.159
R7658 VSS.t2061 VSS.t2007 997.159
R7659 VSS.t4114 VSS.t4098 997.159
R7660 VSS.n715 VSS.t1108 997.159
R7661 VSS.t1328 VSS.t2266 997.159
R7662 VSS.t2371 VSS.t3202 983.311
R7663 VSS.t4317 VSS.t3969 983.311
R7664 VSS.t3549 VSS.t1531 983.311
R7665 VSS.t1325 VSS.t2904 983.311
R7666 VSS.t1557 VSS.t1904 983.311
R7667 VSS.t3314 VSS.t1628 983.311
R7668 VSS.t1809 VSS.t2241 983.311
R7669 VSS.t3471 VSS.t2026 983.311
R7670 VSS.t2305 VSS.t3071 978.693
R7671 VSS.t3138 VSS.t1887 978.693
R7672 VSS.n2429 VSS.n2428 974.801
R7673 VSS.t2369 VSS.t3698 974.077
R7674 VSS.t364 VSS.t1204 969.461
R7675 VSS.t1959 VSS.t331 969.461
R7676 VSS.t4323 VSS.t1320 969.461
R7677 VSS.t1709 VSS.t680 964.845
R7678 VSS.t1276 VSS.t2977 964.845
R7679 VSS.t323 VSS.t3098 964.845
R7680 VSS.t3430 VSS.t1106 964.845
R7681 VSS.t3367 VSS.t4261 964.845
R7682 VSS.t3704 VSS.t3692 964.845
R7683 VSS.n1458 VSS.t2635 955.611
R7684 VSS.t3432 VSS.t1812 946.379
R7685 VSS.t2530 VSS.t2670 946.379
R7686 VSS.t1749 VSS.t0 941.761
R7687 VSS.t692 VSS.t3900 941.761
R7688 VSS.t1116 VSS.t27 941.761
R7689 VSS.t3474 VSS.t26 941.761
R7690 VSS.t652 VSS.t1113 941.761
R7691 VSS.t17 VSS.t851 941.761
R7692 VSS.t2406 VSS.t3700 941.761
R7693 VSS.t757 VSS.t761 941.683
R7694 VSS.t2845 VSS.t3367 937.145
R7695 VSS.t3219 VSS.t1486 937.145
R7696 VSS.t1971 VSS.t796 936.098
R7697 VSS.t501 VSS.t4295 936.098
R7698 VSS.t679 VSS.t3839 932.529
R7699 VSS.t2342 VSS.t38 927.913
R7700 VSS.t2515 VSS.t831 918.679
R7701 VSS.n927 VSS.t1644 918.679
R7702 VSS.n871 VSS.t1037 918.679
R7703 VSS.n800 VSS.t1060 918.679
R7704 VSS.n724 VSS.t3028 918.679
R7705 VSS.n655 VSS.t1938 918.679
R7706 VSS.t1403 VSS.t3049 918.679
R7707 VSS.t3098 VSS.n412 918.679
R7708 VSS.n552 VSS.t3631 918.679
R7709 VSS.t2841 VSS.t36 918.679
R7710 VSS.t2709 VSS.t28 918.679
R7711 VSS.n1516 VSS.t3498 918.679
R7712 VSS.t3514 VSS.n458 918.679
R7713 VSS.t3914 VSS.t3006 918.679
R7714 VSS.t1996 VSS.t501 909.466
R7715 VSS.t2161 VSS.t4087 909.447
R7716 VSS.t1596 VSS.t1126 909.447
R7717 VSS.t3297 VSS.t3635 909.447
R7718 VSS.t491 VSS.t2628 904.831
R7719 VSS.t1124 VSS.t4100 904.831
R7720 VSS.t808 VSS.t2186 904.831
R7721 VSS.t1334 VSS.t484 900.213
R7722 VSS.t3512 VSS.t763 900.213
R7723 VSS.t2980 VSS.t3494 900.213
R7724 VSS.t4259 VSS.t765 900.213
R7725 VSS.t2872 VSS.t849 900.213
R7726 VSS.n2231 VSS.n94 895.597
R7727 VSS.n2424 VSS.n76 895.597
R7728 VSS.n2230 VSS.n359 895.597
R7729 VSS.n2426 VSS.n75 895.597
R7730 VSS.n2229 VSS.n360 895.597
R7731 VSS.n2427 VSS.n74 895.597
R7732 VSS.n2228 VSS.n361 895.597
R7733 VSS.n2429 VSS.n73 895.597
R7734 VSS.n2227 VSS.n362 895.597
R7735 VSS.n2430 VSS.n72 895.597
R7736 VSS.n2226 VSS.n363 895.597
R7737 VSS.t3768 VSS.t1908 895.597
R7738 VSS.n2432 VSS.n71 895.597
R7739 VSS.n2225 VSS.n364 895.597
R7740 VSS.n2434 VSS.n70 895.597
R7741 VSS.n2224 VSS.n365 895.597
R7742 VSS.n2435 VSS.n69 895.597
R7743 VSS.n2223 VSS.n366 895.597
R7744 VSS.n2437 VSS.n68 895.597
R7745 VSS.t18 VSS.t1084 895.597
R7746 VSS.t1121 VSS.t759 895.597
R7747 VSS.n2438 VSS.n67 895.597
R7748 VSS.n2222 VSS.n367 895.597
R7749 VSS.n2440 VSS.n66 895.597
R7750 VSS.n2221 VSS.n368 895.597
R7751 VSS.n2219 VSS.n370 895.597
R7752 VSS.n576 VSS.n575 895.597
R7753 VSS.n579 VSS.n578 895.597
R7754 VSS.n2218 VSS.n371 895.597
R7755 VSS.n2220 VSS.n369 895.597
R7756 VSS.n2133 VSS.n65 895.597
R7757 VSS.t315 VSS.t2272 886.365
R7758 VSS.t321 VSS.t2686 886.365
R7759 VSS.t2472 VSS.t3766 881.747
R7760 VSS.t1966 VSS.t3117 881.747
R7761 VSS.t653 VSS.t2596 881.747
R7762 VSS.t25 VSS.t706 873.801
R7763 VSS.t3096 VSS.t1445 872.514
R7764 VSS.t1743 VSS.t3318 872.514
R7765 VSS.t3720 VSS.t3976 872.514
R7766 VSS.t2034 VSS.t3572 867.899
R7767 VSS.t2544 VSS.t3360 867.899
R7768 VSS.t1307 VSS.t530 867.899
R7769 VSS.t4137 VSS.t2216 867.899
R7770 VSS.t4063 VSS.t299 867.899
R7771 VSS.t167 VSS.t281 867.899
R7772 VSS.t165 VSS.t1332 867.899
R7773 VSS.t2125 VSS.t1124 867.899
R7774 VSS.t813 VSS.t3065 867.899
R7775 VSS.t13 VSS.t1870 867.899
R7776 VSS.t1107 VSS.t648 864.884
R7777 VSS.t2562 VSS.t2375 863.282
R7778 VSS.t3831 VSS.t167 863.282
R7779 VSS.t4158 VSS.t3170 863.282
R7780 VSS.t4188 VSS.t2484 854.048
R7781 VSS.t1969 VSS.t3716 851.51
R7782 VSS.t1692 VSS.t4305 849.433
R7783 VSS.t2223 VSS.t4309 849.433
R7784 VSS.t2387 VSS.t1042 849.433
R7785 VSS.t3655 VSS.t1050 849.433
R7786 VSS.t3786 VSS.t1054 849.433
R7787 VSS.t1694 VSS.t1046 849.433
R7788 VSS.t3200 VSS.n1716 849.433
R7789 VSS.t2611 VSS.t4184 849.433
R7790 VSS.n1717 VSS.t3791 849.433
R7791 VSS.t544 VSS.t3040 849.433
R7792 VSS.t3198 VSS.t2035 849.433
R7793 VSS.t2315 VSS.t4195 849.433
R7794 VSS.t1272 VSS.t1990 849.433
R7795 VSS.t283 VSS.t2005 849.433
R7796 VSS.t1910 VSS.t3684 849.433
R7797 VSS.n1851 VSS.t2678 849.433
R7798 VSS.t840 VSS.n1851 849.433
R7799 VSS.t1908 VSS.t1859 849.433
R7800 VSS.t5 VSS.t958 849.433
R7801 VSS.t425 VSS.t467 849.433
R7802 VSS.t1130 VSS.t839 849.433
R7803 VSS.t1858 VSS.t4188 849.433
R7804 VSS.t3900 VSS.t3945 849.433
R7805 VSS.t2173 VSS.t3584 849.433
R7806 VSS.n800 VSS.t2361 849.433
R7807 VSS.t1108 VSS.t1098 849.433
R7808 VSS.t1096 VSS.t1115 849.433
R7809 VSS.n724 VSS.t1967 849.433
R7810 VSS.t994 VSS.t3183 849.433
R7811 VSS.t658 VSS.n708 849.433
R7812 VSS.t1081 VSS.t23 849.433
R7813 VSS.t3104 VSS.t3899 849.433
R7814 VSS.t3565 VSS.t1889 849.433
R7815 VSS.t3696 VSS.t837 849.433
R7816 VSS.t325 VSS.n412 849.433
R7817 VSS.t392 VSS.n419 849.433
R7818 VSS.t4200 VSS.n399 849.433
R7819 VSS.t654 VSS.t3306 849.433
R7820 VSS.n458 VSS.t406 849.433
R7821 VSS.t1660 VSS.t3876 849.433
R7822 VSS.t2025 VSS.t2303 844.816
R7823 VSS.n576 VSS.n65 843.15
R7824 VSS.n980 VSS.t533 835.582
R7825 VSS.t4195 VSS.t2544 835.582
R7826 VSS.t3738 VSS.t3348 835.582
R7827 VSS.t3316 VSS.t2845 835.582
R7828 VSS.t4267 VSS.t691 830.966
R7829 VSS.t2655 VSS.t526 830.966
R7830 VSS.t3669 VSS.t4061 830.966
R7831 VSS.t3557 VSS.t688 830.966
R7832 VSS.t1 VSS.t311 830.966
R7833 VSS.t2274 VSS.t309 830.966
R7834 VSS.t1625 VSS.t315 830.966
R7835 VSS.t2649 VSS.t425 830.966
R7836 VSS.t1222 VSS.t3756 830.966
R7837 VSS.t493 VSS.t159 830.966
R7838 VSS.t4194 VSS.t147 830.966
R7839 VSS.t812 VSS.t149 830.966
R7840 VSS.t2690 VSS.t678 830.966
R7841 VSS.t2988 VSS.t3045 830.966
R7842 VSS.t1527 VSS.t500 830.966
R7843 VSS.t3744 VSS.t3008 830.966
R7844 VSS.t179 VSS.t963 830.966
R7845 VSS.t1640 VSS.t792 830.966
R7846 VSS.t1147 VSS.t3475 830.966
R7847 VSS.t844 VSS.t2394 826.35
R7848 VSS.t2470 VSS.t1130 826.35
R7849 VSS.t24 VSS.t1082 820.303
R7850 VSS.t3028 VSS.t1966 817.116
R7851 VSS.t2596 VSS.t1077 817.116
R7852 VSS.t1594 VSS.t653 817.116
R7853 VSS.t1413 VSS.t3461 817.116
R7854 VSS.t3702 VSS.t1572 817.116
R7855 VSS.t1514 VSS.t4057 812.5
R7856 VSS.t366 VSS.n865 812.5
R7857 VSS.t16 VSS.t1111 812.5
R7858 VSS.t3686 VSS.t3897 807.885
R7859 VSS.t2746 VSS.t4294 807.885
R7860 VSS.t1948 VSS.t4007 803.268
R7861 VSS.t3899 VSS.t4182 803.268
R7862 VSS.t126 VSS.t1528 798.652
R7863 VSS.t1621 VSS.t1641 798.652
R7864 VSS.t2051 VSS.t690 794.034
R7865 VSS.n1464 VSS.t4091 794.034
R7866 VSS.t1416 VSS.t1862 794.034
R7867 VSS.t1877 VSS.t469 789.418
R7868 VSS.t3516 VSS.t8 789.418
R7869 VSS.n2436 VSS.n2435 785.034
R7870 VSS.t2270 VSS.t793 784.802
R7871 VSS.n2437 VSS.n2436 781.039
R7872 VSS.t4235 VSS.t1509 780.186
R7873 VSS.t3599 VSS.t1091 780.186
R7874 VSS.t1657 VSS.t1655 775.568
R7875 VSS.t3999 VSS.t1408 775.568
R7876 VSS.t530 VSS.t2519 775.568
R7877 VSS.t487 VSS.t3614 775.568
R7878 VSS.t932 VSS.t933 775.568
R7879 VSS.t4359 VSS.t4361 775.568
R7880 VSS.t1267 VSS.t1269 775.568
R7881 VSS.t2641 VSS.t2643 775.568
R7882 VSS.t527 VSS.t3928 775.568
R7883 VSS.t3928 VSS.t3926 775.568
R7884 VSS.t3156 VSS.t3155 775.568
R7885 VSS.t1518 VSS.t3669 775.568
R7886 VSS.t2154 VSS.t779 775.568
R7887 VSS.t3823 VSS.t2154 775.568
R7888 VSS.t2715 VSS.t2713 775.568
R7889 VSS.t2291 VSS.t2290 775.568
R7890 VSS.t3377 VSS.t3375 775.568
R7891 VSS.t1815 VSS.t1816 775.568
R7892 VSS.t3542 VSS.t3540 775.568
R7893 VSS.t2310 VSS.t2309 775.568
R7894 VSS.t3941 VSS.t3943 775.568
R7895 VSS.t478 VSS.t1168 775.568
R7896 VSS.t3609 VSS.t3607 775.568
R7897 VSS.t549 VSS.t3266 775.568
R7898 VSS.t2826 VSS.t141 775.568
R7899 VSS.t2199 VSS.t489 775.568
R7900 VSS.t987 VSS.t988 775.568
R7901 VSS.t547 VSS.t2215 775.568
R7902 VSS.t1452 VSS.t1454 775.568
R7903 VSS.t551 VSS.t3079 775.568
R7904 VSS.t1193 VSS.t1191 775.568
R7905 VSS.t3473 VSS.t137 775.568
R7906 VSS.t3472 VSS.t135 775.568
R7907 VSS.t2647 VSS.t1702 775.568
R7908 VSS.t2646 VSS.t2647 775.568
R7909 VSS.t3568 VSS.t3570 775.568
R7910 VSS.t1389 VSS.t3568 775.568
R7911 VSS.t517 VSS.t3410 775.568
R7912 VSS.t2775 VSS.t2948 775.568
R7913 VSS.t2606 VSS.t777 775.568
R7914 VSS.t829 VSS.t3169 775.568
R7915 VSS.t1317 VSS.t1315 775.568
R7916 VSS.t1799 VSS.t1800 775.568
R7917 VSS.t2023 VSS.t2025 775.568
R7918 VSS.t775 VSS.t2859 775.568
R7919 VSS.t2859 VSS.t4092 775.568
R7920 VSS.t1449 VSS.t1451 775.568
R7921 VSS.t1007 VSS.t1999 775.568
R7922 VSS.t773 VSS.t919 775.568
R7923 VSS.t3193 VSS.t3194 775.568
R7924 VSS.t3276 VSS.t3278 775.568
R7925 VSS.t553 VSS.t2954 775.568
R7926 VSS.t1929 VSS.t1927 775.568
R7927 VSS.t797 VSS.t4097 775.568
R7928 VSS.t4097 VSS.t2822 775.568
R7929 VSS.t801 VSS.t3301 775.568
R7930 VSS.t781 VSS.t1466 775.568
R7931 VSS.t2177 VSS.t2178 775.568
R7932 VSS.t3530 VSS.t3532 775.568
R7933 VSS.t3127 VSS.t3128 775.568
R7934 VSS.t4315 VSS.t4313 775.568
R7935 VSS.t1486 VSS.t2580 775.568
R7936 VSS.t2839 VSS.t2838 775.568
R7937 VSS.t2823 VSS.t2824 775.568
R7938 VSS.t785 VSS.t1517 775.568
R7939 VSS.t1542 VSS.t1541 775.568
R7940 VSS.t3862 VSS.t3864 775.568
R7941 VSS.t2581 VSS.t2582 775.568
R7942 VSS.t4294 VSS.t4292 775.568
R7943 VSS.t2612 VSS.t1229 770.952
R7944 VSS.t2502 VSS.t4106 770.952
R7945 VSS.t1686 VSS.t2014 770.952
R7946 VSS.t2206 VSS.t2488 770.952
R7947 VSS.t128 VSS.t3545 770.952
R7948 VSS.t1085 VSS.t3822 766.336
R7949 VSS.t3777 VSS.t502 761.72
R7950 VSS.t2352 VSS.t537 761.72
R7951 VSS.t1100 VSS.t3718 757.102
R7952 VSS.t1094 VSS.t755 757.102
R7953 VSS.t1098 VSS.t751 757.102
R7954 VSS.t1517 VSS.n614 757.102
R7955 VSS.t504 VSS.t2310 747.87
R7956 VSS.t1967 VSS.t3836 747.87
R7957 VSS.t1702 VSS.t2914 747.87
R7958 VSS.t815 VSS.t3221 747.386
R7959 VSS.t2748 VSS.t539 747.386
R7960 VSS.t3269 VSS.t4089 743.254
R7961 VSS.t2824 VSS.t4235 743.254
R7962 VSS.t469 VSS.n794 738.636
R7963 VSS.t1970 VSS.t3496 738.636
R7964 VSS.t918 VSS.t3490 738.636
R7965 VSS.t1636 VSS.t3492 738.636
R7966 VSS.t2888 VSS.t2680 734.02
R7967 VSS.t680 VSS.t2579 734.02
R7968 VSS.t2450 VSS.t323 734.02
R7969 VSS.t1106 VSS.t1407 734.02
R7970 VSS.t4261 VSS.t1228 734.02
R7971 VSS.t856 VSS.t850 731.139
R7972 VSS.t858 VSS.t857 731.139
R7973 VSS.t2451 VSS.t1997 731.139
R7974 VSS.t1105 VSS.t1119 729.404
R7975 VSS.t657 VSS.t647 729.404
R7976 VSS.t3071 VSS.t673 724.788
R7977 VSS.t1159 VSS.t2662 724.788
R7978 VSS.t4007 VSS.n648 724.788
R7979 VSS.t480 VSS.t1447 724.788
R7980 VSS.t3815 VSS.t1513 720.17
R7981 VSS.t3809 VSS.t2109 720.17
R7982 VSS.t3811 VSS.t3387 720.17
R7983 VSS.t232 VSS.t3558 720.17
R7984 VSS.t2316 VSS.t1751 720.17
R7985 VSS.t1751 VSS.t509 720.17
R7986 VSS.t430 VSS.t3866 720.17
R7987 VSS.t432 VSS.t4030 720.17
R7988 VSS.t428 VSS.t2996 720.17
R7989 VSS.t4215 VSS.t3152 720.17
R7990 VSS.t3574 VSS.t3578 720.17
R7991 VSS.t2590 VSS.t1584 720.17
R7992 VSS.t3774 VSS.t885 720.17
R7993 VSS.t909 VSS.t3351 720.17
R7994 VSS.t607 VSS.t1805 720.17
R7995 VSS.t907 VSS.t1066 720.17
R7996 VSS.t3640 VSS.t1865 720.17
R7997 VSS.t777 VSS.t3640 720.17
R7998 VSS.t3421 VSS.t829 720.17
R7999 VSS.t3034 VSS.t3421 720.17
R8000 VSS.t1680 VSS.t3439 720.17
R8001 VSS.t1672 VSS.t3434 720.17
R8002 VSS.t1676 VSS.t3784 720.17
R8003 VSS.t177 VSS.t2550 720.17
R8004 VSS.t181 VSS.t1008 720.17
R8005 VSS.t185 VSS.t3299 720.17
R8006 VSS.t3653 VSS.t4014 720.17
R8007 VSS.t4014 VSS.t821 720.17
R8008 VSS.t3603 VSS.t4218 720.17
R8009 VSS.t673 VSS.t498 715.554
R8010 VSS.t2129 VSS.t4317 715.554
R8011 VSS.t2874 VSS.t2880 715.554
R8012 VSS.t1946 VSS.t2031 715.554
R8013 VSS.t362 VSS.t1202 710.938
R8014 VSS.t1961 VSS.t368 710.938
R8015 VSS.t1620 VSS.t3214 706.322
R8016 VSS.t1618 VSS.t3212 706.322
R8017 VSS.t2864 VSS.t1193 706.322
R8018 VSS.t2008 VSS.t1317 706.322
R8019 VSS.t4334 VSS.t685 701.706
R8020 VSS.t4008 VSS.t4187 701.706
R8021 VSS.t996 VSS.t367 701.706
R8022 VSS.t2260 VSS.t4197 701.706
R8023 VSS.t525 VSS.t2385 701.706
R8024 VSS.t1644 VSS.t1944 701.706
R8025 VSS.t1037 VSS.t2061 701.706
R8026 VSS.t4186 VSS.t1479 701.706
R8027 VSS.n794 VSS.t2601 701.706
R8028 VSS.t1895 VSS.t1149 701.706
R8029 VSS.t1012 VSS.t3868 701.706
R8030 VSS.t2075 VSS.t4075 701.706
R8031 VSS.t873 VSS.t1116 701.706
R8032 VSS.t924 VSS.t2722 701.706
R8033 VSS.t1009 VSS.n390 701.706
R8034 VSS.t1070 VSS.n622 701.706
R8035 VSS.t3075 VSS.t3565 697.088
R8036 VSS.t2805 VSS.t42 697.088
R8037 VSS.t1083 VSS.t704 695.473
R8038 VSS.n905 VSS.t3269 692.472
R8039 VSS.t2532 VSS.t2666 687.856
R8040 VSS.t1383 VSS.t4220 687.856
R8041 VSS.t3674 VSS.t514 683.24
R8042 VSS.t2558 VSS.t4133 683.24
R8043 VSS.t293 VSS.t1860 683.24
R8044 VSS.t1331 VSS.t2044 683.24
R8045 VSS.t877 VSS.t869 683.24
R8046 VSS.t881 VSS.t859 683.24
R8047 VSS.t875 VSS.t861 683.24
R8048 VSS.t1285 VSS.t835 683.24
R8049 VSS.t1153 VSS.t4079 683.24
R8050 VSS.t2890 VSS.t3042 678.622
R8051 VSS.t4192 VSS.t171 678.622
R8052 VSS.t4162 VSS.t1073 678.622
R8053 VSS.t767 VSS.t1079 678.622
R8054 VSS.t1900 VSS.t799 678.622
R8055 VSS.t1324 VSS.t1085 674.006
R8056 VSS.t3573 VSS.t1982 669.389
R8057 VSS.t3668 VSS.t2502 669.389
R8058 VSS.t3365 VSS.t2243 669.389
R8059 VSS.t1889 VSS.t770 669.389
R8060 VSS.t2106 VSS.t1604 664.774
R8061 VSS.t2688 VSS.t1598 664.774
R8062 VSS.t2217 VSS.t3724 664.774
R8063 VSS.t681 VSS.t4223 664.774
R8064 VSS.t4285 VSS.t470 664.774
R8065 VSS.t3447 VSS.t2813 664.774
R8066 VSS.t4032 VSS.t52 664.774
R8067 VSS.t702 VSS.t684 664.774
R8068 VSS.t665 VSS.t1118 664.774
R8069 VSS.t131 VSS.t3055 664.774
R8070 VSS.t1803 VSS.t911 664.774
R8071 VSS.t2948 VSS.t3420 664.774
R8072 VSS.t3371 VSS.t800 664.774
R8073 VSS.t1525 VSS.t832 664.774
R8074 VSS.t3436 VSS.t1674 664.774
R8075 VSS.t475 VSS.t916 664.774
R8076 VSS.t663 VSS.t400 664.774
R8077 VSS.t1868 VSS.t4202 664.774
R8078 VSS.t4198 VSS.t1009 664.774
R8079 VSS.t1642 VSS.t803 664.774
R8080 VSS.t3107 VSS.t2124 664.774
R8081 VSS.t1574 VSS.t2975 664.774
R8082 VSS.t3404 VSS.t1128 664.774
R8083 VSS.t1402 VSS.t1932 660.157
R8084 VSS.t2609 VSS.t2298 660.157
R8085 VSS.t2708 VSS.t30 660.157
R8086 VSS.t3155 VSS.t2910 655.54
R8087 VSS.t1630 VSS.t2221 655.54
R8088 VSS.t3308 VSS.t535 655.54
R8089 VSS.t1888 VSS.t4245 650.923
R8090 VSS.t3631 VSS.t1980 650.923
R8091 VSS.t690 VSS.t4000 646.308
R8092 VSS.n1464 VSS.t3061 646.308
R8093 VSS.t1570 VSS.t3082 641.691
R8094 VSS.t2127 VSS.t2537 641.691
R8095 VSS.t467 VSS.t4034 641.691
R8096 VSS.t3898 VSS.t2280 641.691
R8097 VSS.t1792 VSS.t2029 641.691
R8098 VSS.n577 VSS.n576 640.429
R8099 VSS.t3685 VSS.t2627 637.074
R8100 VSS.n1852 VSS.t3768 632.457
R8101 VSS.t3498 VSS.t3283 632.457
R8102 VSS.t3847 VSS.t3795 632.457
R8103 VSS.t4057 VSS.t1004 627.841
R8104 VSS.t3830 VSS.t1280 618.609
R8105 VSS.t3128 VSS.t1041 618.609
R8106 VSS.t2394 VSS.t366 613.991
R8107 VSS.t4049 VSS.t3758 613.991
R8108 VSS.t1072 VSS.t4040 613.991
R8109 VSS.t2635 VSS.t3297 613.991
R8110 VSS.t3865 VSS.t1222 609.375
R8111 VSS.t3352 VSS.t2988 609.375
R8112 VSS.t3438 VSS.t3744 609.375
R8113 VSS.t3300 VSS.t179 609.375
R8114 VSS.t2560 VSS.t2365 604.76
R8115 VSS.t2396 VSS.t4074 604.76
R8116 VSS.t422 VSS.t3667 604.76
R8117 VSS.t3348 VSS.t1006 604.76
R8118 VSS.t3399 VSS.t545 604.76
R8119 VSS.t38 VSS.t2806 595.527
R8120 VSS.t3597 VSS.t833 595.527
R8121 VSS.n2428 VSS.n2427 591.273
R8122 VSS.t4000 VSS.t3198 590.909
R8123 VSS.t27 VSS.t139 590.909
R8124 VSS.t2738 VSS.t2301 590.909
R8125 VSS.t1912 VSS.t1187 586.293
R8126 VSS.t1191 VSS.t2567 586.293
R8127 VSS.t1800 VSS.t3415 586.293
R8128 VSS.t3700 VSS.t3527 581.677
R8129 VSS.t3306 VSS.t1158 577.061
R8130 VSS.t2152 VSS.t932 577.061
R8131 VSS.t1812 VSS.t4359 577.061
R8132 VSS.t2670 VSS.t2950 577.061
R8133 VSS.t3162 VSS.t1007 577.061
R8134 VSS.t3340 VSS.t3847 577.061
R8135 VSS.t1004 VSS.t1307 572.443
R8136 VSS.t2617 VSS.t317 572.443
R8137 VSS.t2215 VSS.t3328 572.443
R8138 VSS.t1157 VSS.t3594 572.443
R8139 VSS.t2660 VSS.t1160 567.827
R8140 VSS.t3010 VSS.t4042 567.827
R8141 VSS.t998 VSS.t2839 567.827
R8142 VSS.t3196 VSS.t1023 567.827
R8143 VSS.t2498 VSS.t2279 567.827
R8144 VSS.t533 VSS.t3685 563.211
R8145 VSS.n2441 VSS.n65 559.232
R8146 VSS.t850 VSS.t854 559.059
R8147 VSS.t3579 VSS.t994 558.595
R8148 VSS.t1122 VSS.t823 558.595
R8149 VSS.t3976 VSS.t2480 558.595
R8150 VSS.t3828 VSS.t2678 553.977
R8151 VSS.t1092 VSS.t747 553.977
R8152 VSS.t3570 VSS.t2646 553.977
R8153 VSS.t2776 VSS.t21 553.977
R8154 VSS.t3419 VSS.t3643 553.977
R8155 VSS.t2860 VSS.t2878 553.977
R8156 VSS.t1385 VSS.t2012 553.977
R8157 VSS.t838 VSS.t3849 549.361
R8158 VSS.n1995 VSS.t2476 549.361
R8159 VSS.t2087 VSS.t3308 544.745
R8160 VSS.t2630 VSS.t1554 540.129
R8161 VSS.t988 VSS.t1557 540.129
R8162 VSS.t2188 VSS.t1867 540.129
R8163 VSS.t1927 VSS.t1809 540.129
R8164 VSS.t2597 VSS.t1729 535.511
R8165 VSS.t2959 VSS.t1717 535.511
R8166 VSS.t3175 VSS.t1725 535.511
R8167 VSS.t4273 VSS.t1723 535.511
R8168 VSS.t1234 VSS.t4267 535.511
R8169 VSS.t3789 VSS.t2489 535.511
R8170 VSS.t1646 VSS.t1248 535.511
R8171 VSS.t842 VSS.t1324 535.511
R8172 VSS.t1035 VSS.t2002 535.511
R8173 VSS.n1333 VSS.t4158 535.511
R8174 VSS.t2122 VSS.t855 535.511
R8175 VSS.t3420 VSS.t1205 535.511
R8176 VSS.t2589 VSS.t1411 535.511
R8177 VSS.t1696 VSS.t3112 535.511
R8178 VSS.t511 VSS.t3573 530.895
R8179 VSS.t2921 VSS.t3168 526.279
R8180 VSS.n2423 VSS.t626 522.259
R8181 VSS.n2425 VSS.t89 522.259
R8182 VSS.n2428 VSS.t1368 522.259
R8183 VSS.n2431 VSS.t1844 522.259
R8184 VSS.n2433 VSS.t240 522.259
R8185 VSS.n2439 VSS.t573 522.259
R8186 VSS.n2436 VSS.t739 522.259
R8187 VSS.n2444 VSS.t728 522.259
R8188 VSS.n2448 VSS.t1835 522.259
R8189 VSS.n2452 VSS.t80 522.259
R8190 VSS.n2454 VSS.t617 522.259
R8191 VSS.n2450 VSS.t1359 522.259
R8192 VSS.n2446 VSS.t261 522.259
R8193 VSS.n2442 VSS.t599 522.259
R8194 VSS.t519 VSS.t1576 521.663
R8195 VSS.t3901 VSS.t863 521.663
R8196 VSS.t2838 VSS.t2496 521.663
R8197 VSS.n2426 VSS.n2425 517.364
R8198 VSS.t2927 VSS.t3888 517.045
R8199 VSS.t3904 VSS.t977 517.045
R8200 VSS.t1973 VSS.t1698 517.045
R8201 VSS.t3036 VSS.t3476 517.045
R8202 VSS.t3147 VSS.t2651 517.045
R8203 VSS.t2884 VSS.t3970 517.045
R8204 VSS.t4001 VSS.t2454 517.045
R8205 VSS.t2040 VSS.t3974 517.045
R8206 VSS.t4328 VSS.t3510 517.045
R8207 VSS.t3355 VSS.t1238 517.045
R8208 VSS.t1246 VSS.t3895 517.045
R8209 VSS.t3872 VSS.t2391 517.045
R8210 VSS.t3525 VSS.t4340 517.045
R8211 VSS.t2057 VSS.t2524 517.045
R8212 VSS.t1183 VSS.t1342 517.045
R8213 VSS.t2379 VSS.t2059 517.045
R8214 VSS.t1707 VSS.t1185 517.045
R8215 VSS.t1653 VSS.t2293 517.045
R8216 VSS.t2110 VSS.t3206 517.045
R8217 VSS.t2276 VSS.t3444 517.045
R8218 VSS.t3149 VSS.t3249 517.045
R8219 VSS.t1293 VSS.t1495 517.045
R8220 VSS.t2032 VSS.t1873 517.045
R8221 VSS.t1289 VSS.t3906 517.045
R8222 VSS.t2167 VSS.t3245 517.045
R8223 VSS.t3563 VSS.t1300 517.045
R8224 VSS.t1505 VSS.t3860 517.045
R8225 VSS.t3953 VSS.t4124 517.045
R8226 VSS.t3408 VSS.t928 517.045
R8227 VSS.t2886 VSS.t3854 517.045
R8228 VSS.t1757 VSS.t2504 517.045
R8229 VSS.t2548 VSS.t1460 517.045
R8230 VSS.t1419 VSS.t3402 517.045
R8231 VSS.t3426 VSS.t2246 517.045
R8232 VSS.t3231 VSS.t1236 517.045
R8233 VSS.t1232 VSS.t2139 517.045
R8234 VSS.t2552 VSS.t1464 517.045
R8235 VSS.t3255 VSS.t2491 517.045
R8236 VSS.t3087 VSS.t3972 517.045
R8237 VSS.t1533 VSS.t4128 517.045
R8238 VSS.t2999 VSS.t1992 517.045
R8239 VSS.t3210 VSS.t1029 517.045
R8240 VSS.t3752 VSS.t3566 517.045
R8241 VSS.t965 VSS.t3229 517.045
R8242 VSS.t2535 VSS.t3166 517.045
R8243 VSS.t973 VSS.t3122 517.045
R8244 VSS.t2180 VSS.t1392 517.045
R8245 VSS.t1529 VSS.t3486 517.045
R8246 VSS.t3694 VSS.t3886 517.045
R8247 VSS.t2898 VSS.t3726 517.045
R8248 VSS.t1212 VSS.t4231 517.045
R8249 VSS.t3100 VSS.t1261 517.045
R8250 VSS.t3949 VSS.t1278 517.045
R8251 VSS.t4321 VSS.t3189 517.045
R8252 VSS.t4251 VSS.t2906 517.045
R8253 VSS.t1139 VSS.t3032 517.045
R8254 VSS.t1473 VSS.t985 517.045
R8255 VSS.t954 VSS.t1638 517.045
R8256 VSS.t2468 VSS.t2957 517.045
R8257 VSS.t1000 VSS.t1987 517.045
R8258 VSS.t1291 VSS.t2322 517.045
R8259 VSS.t2233 VSS.t1387 517.045
R8260 VSS.t2493 VSS.t1295 517.045
R8261 VSS.t2900 VSS.t2286 517.045
R8262 VSS.t3038 VSS.t1983 517.045
R8263 VSS.t4216 VSS.t2827 517.045
R8264 VSS.t1634 VSS.t3457 517.045
R8265 VSS.t3451 VSS.t2770 517.045
R8266 VSS.t2159 VSS.t2657 517.045
R8267 VSS.t4018 VSS.t1586 517.045
R8268 VSS.t2604 VSS.t2965 517.045
R8269 VSS.t2973 VSS.t3935 517.045
R8270 VSS.t3924 VSS.t2016 517.045
R8271 VSS.t956 VSS.t1715 517.045
R8272 VSS.t3488 VSS.t3251 517.045
R8273 VSS.t2607 VSS.t3285 517.045
R8274 VSS.t2694 VSS.t3931 517.045
R8275 VSS.t2835 VSS.t1151 517.045
R8276 VSS.t1477 VSS.t2353 517.045
R8277 VSS.t3891 VSS.t2284 517.045
R8278 VSS.t2952 VSS.t2554 517.045
R8279 VSS.t3625 VSS.t2163 517.045
R8280 VSS.t3464 VSS.t2961 517.045
R8281 VSS.t3762 VSS.t2466 517.045
R8282 VSS.t1177 VSS.t2346 517.045
R8283 VSS.t992 VSS.t2633 517.045
R8284 VSS.t541 VSS.t4139 517.045
R8285 VSS.t3550 VSS.t2081 517.045
R8286 VSS.t2526 VSS.t2288 517.045
R8287 VSS.t2182 VSS.t1755 517.045
R8288 VSS.t3627 VSS.t3389 517.045
R8289 VSS.t2211 VSS.t1143 517.045
R8290 VSS.t3118 VSS.t4151 517.045
R8291 VSS.t4275 VSS.t2772 517.045
R8292 VSS.t3334 VSS.t3963 517.045
R8293 VSS.t1852 VSS.t1918 517.045
R8294 VSS.t1336 VSS.t4176 517.045
R8295 VSS.t3018 VSS.t2063 517.045
R8296 VSS.t1251 VSS.t1770 517.045
R8297 VSS.t3338 VSS.t1405 517.045
R8298 VSS.t2131 VSS.t3083 517.045
R8299 VSS.t1226 VSS.t3712 517.045
R8300 VSS.t3233 VSS.t2711 517.045
R8301 VSS.t2069 VSS.t2042 517.045
R8302 VSS.t2118 VSS.t1763 517.045
R8303 VSS.t4241 VSS.t3073 517.045
R8304 VSS.t1021 VSS.t2963 517.045
R8305 VSS.t3561 VSS.t1807 517.045
R8306 VSS.t4355 VSS.t2785 517.045
R8307 VSS.t1374 VSS.t2938 517.045
R8308 VSS.t2594 VSS.t1033 517.045
R8309 VSS.t3241 VSS.t4122 517.045
R8310 VSS.t3484 VSS.t2462 517.045
R8311 VSS.t1458 VSS.t1940 517.045
R8312 VSS.t3519 VSS.t1914 517.045
R8313 VSS.t3440 VSS.t1772 517.045
R8314 VSS.t3181 VSS.t2478 517.045
R8315 VSS.t2328 VSS.t4077 517.045
R8316 VSS.t1958 VSS.t4135 517.045
R8317 VSS.t3791 VSS.t1377 517.045
R8318 VSS.t2894 VSS.t3125 517.045
R8319 VSS.t2720 VSS.t3554 517.045
R8320 VSS.t4350 VSS.t2235 517.045
R8321 VSS.t2971 VSS.t2448 517.045
R8322 VSS.t3067 VSS.t1214 517.045
R8323 VSS.t2870 VSS.t3047 517.045
R8324 VSS.t2724 VSS.t3191 517.045
R8325 VSS.t4239 VSS.t3324 517.045
R8326 VSS.t952 VSS.t2146 517.045
R8327 VSS.t3521 VSS.t1774 517.045
R8328 VSS.t3649 VSS.t3916 517.045
R8329 VSS.t2702 VSS.t3417 517.045
R8330 VSS.t1002 VSS.t3411 517.045
R8331 VSS.t1297 VSS.t1881 517.045
R8332 VSS.t2258 VSS.t2969 517.045
R8333 VSS.t2934 VSS.t1421 517.045
R8334 VSS.t4297 VSS.t1253 517.045
R8335 VSS.t3740 VSS.t3714 517.045
R8336 VSS.t3793 VSS.t3615 517.045
R8337 VSS.t3077 VSS.t3462 517.045
R8338 VSS.t2540 VSS.t3672 517.045
R8339 VSS.t3094 VSS.t2696 517.045
R8340 VSS.t1244 VSS.t2508 517.045
R8341 VSS.t1507 VSS.n972 517.045
R8342 VSS.t1590 VSS.t3502 517.045
R8343 VSS.t1515 VSS.t4283 517.045
R8344 VSS.t4005 VSS.t3508 517.045
R8345 VSS.t1031 VSS.t2866 517.045
R8346 VSS.t2622 VSS.t1614 517.045
R8347 VSS.t3750 VSS.t960 517.045
R8348 VSS.t1651 VSS.t4287 517.045
R8349 VSS.t2202 VSS.t1705 517.045
R8350 VSS.t3664 VSS.t3043 517.045
R8351 VSS.t2200 VSS.t2510 517.045
R8352 VSS.t3623 VSS.t1481 517.045
R8353 VSS.t1548 VSS.t1608 517.045
R8354 VSS.t3533 VSS.t3644 517.045
R8355 VSS.t3841 VSS.t3243 517.045
R8356 VSS.t2631 VSS.t2165 517.045
R8357 VSS.t2282 VSS.t1883 517.045
R8358 VSS.t979 VSS.t4051 517.045
R8359 VSS.t1964 VSS.t2546 517.045
R8360 VSS.t3177 VSS.t3834 517.045
R8361 VSS.t2157 VSS.t2018 517.045
R8362 VSS.t3145 VSS.t3552 517.045
R8363 VSS.t1027 VSS.t1588 517.045
R8364 VSS.t3311 VSS.t4120 517.045
R8365 VSS.t3678 VSS.t3059 517.045
R8366 VSS.t1179 VSS.t1759 517.045
R8367 VSS.t3153 VSS.t2803 517.045
R8368 VSS.t3619 VSS.t3506 517.045
R8369 VSS.t4243 VSS.t3272 517.045
R8370 VSS.t3582 VSS.t2728 517.045
R8371 VSS.t3024 VSS.t1200 517.045
R8372 VSS.t4022 VSS.t3014 517.045
R8373 VSS.t3393 VSS.t2698 517.045
R8374 VSS.t2908 VSS.t2730 517.045
R8375 VSS.t1662 VSS.t4028 517.045
R8376 VSS.t4069 VSS.t4016 517.045
R8377 VSS.t3884 VSS.t4172 517.045
R8378 VSS.t3710 VSS.t2569 517.045
R8379 VSS.t3326 VSS.t3764 517.045
R8380 VSS.t2350 VSS.t3850 517.045
R8381 VSS.t2833 VSS.t4301 517.045
R8382 VSS.t3459 VSS.t2783 517.045
R8383 VSS.t2936 VSS.t2389 517.045
R8384 VSS.t2359 VSS.t3235 517.045
R8385 VSS.t2777 VSS.t2148 517.045
R8386 VSS.t4093 VSS.t2851 517.045
R8387 VSS.t4010 VSS.t2902 517.045
R8388 VSS.t2102 VSS.t975 517.045
R8389 VSS.t4225 VSS.t3621 517.045
R8390 VSS.t3621 VSS.t4140 517.045
R8391 VSS.t2613 VSS.t3682 517.045
R8392 VSS.t2916 VSS.t3658 517.045
R8393 VSS.t2918 VSS.t3657 517.045
R8394 VSS.t3261 VSS.t2020 517.045
R8395 VSS.t3259 VSS.t2021 517.045
R8396 VSS.t1462 VSS.t3259 517.045
R8397 VSS.t4303 VSS.t1462 517.045
R8398 VSS.t3817 VSS.t3397 517.045
R8399 VSS.t2882 VSS.t3937 517.045
R8400 VSS.t2932 VSS.t1396 517.045
R8401 VSS.t1145 VSS.t4344 517.045
R8402 VSS.t1648 VSS.t1544 517.045
R8403 VSS.t3353 VSS.t3227 517.045
R8404 VSS.t3223 VSS.t2857 517.045
R8405 VSS.t3617 VSS.t3160 517.045
R8406 VSS.t2736 VSS.t1713 517.045
R8407 VSS.t3237 VSS.t2330 517.045
R8408 VSS.t1916 VSS.t2332 517.045
R8409 VSS.t3089 VSS.t1539 517.045
R8410 VSS.t1467 VSS.t3302 517.045
R8411 VSS.t2718 VSS.t1281 517.045
R8412 VSS.t3826 VSS.t3363 517.045
R8413 VSS.t1885 VSS.t2204 517.045
R8414 VSS.t3660 VSS.t2615 517.045
R8415 VSS.t3922 VSS.t3722 517.045
R8416 VSS.t2175 VSS.t3349 517.045
R8417 VSS.t3102 VSS.t3965 517.045
R8418 VSS.t4067 VSS.t4271 517.045
R8419 VSS.t3304 VSS.t3468 517.045
R8420 VSS.t1893 VSS.t2876 517.045
R8421 VSS.t3832 VSS.t2592 517.045
R8422 VSS.t2197 VSS.t2381 517.045
R8423 VSS.t2100 VSS.t4332 517.045
R8424 VSS.t4279 VSS.t3423 517.045
R8425 VSS.t3413 VSS.t3142 517.045
R8426 VSS.t1338 VSS.t3535 517.045
R8427 VSS.t3662 VSS.t1469 517.045
R8428 VSS.t2418 VSS.t1499 517.045
R8429 VSS.t3085 VSS.t1930 517.045
R8430 VSS.t4257 VSS.t3264 517.045
R8431 VSS.t3185 VSS.t2446 517.045
R8432 VSS.t1326 VSS.t4178 517.045
R8433 VSS.t2456 VSS.t3601 517.045
R8434 VSS.t3225 VSS.t1920 517.045
R8435 VSS.t4145 VSS.t3893 517.045
R8436 VSS.t2726 VSS.t3730 517.045
R8437 VSS.t2896 VSS.t2625 517.045
R8438 VSS.t2940 VSS.t3880 517.045
R8439 VSS.t4149 VSS.t1409 517.045
R8440 VSS.t1136 VSS.t1616 517.045
R8441 VSS.t2704 VSS.t1666 517.045
R8442 VSS.t1283 VSS.t2644 517.045
R8443 VSS.t4143 VSS.t3391 517.045
R8444 VSS.t1950 VSS.t293 517.045
R8445 VSS.t305 VSS.t1950 517.045
R8446 VSS.t2189 VSS.t1379 517.045
R8447 VSS.t2945 VSS.t2189 517.045
R8448 VSS.t1014 VSS.t2945 517.045
R8449 VSS.t1016 VSS.t2947 517.045
R8450 VSS.t3001 VSS.t1024 517.045
R8451 VSS.t3002 VSS.t1025 517.045
R8452 VSS.t1501 VSS.t3004 517.045
R8453 VSS.t2239 VSS.t4353 517.045
R8454 VSS.t2984 VSS.t2892 517.045
R8455 VSS.t2104 VSS.t4338 517.045
R8456 VSS.t1394 VSS.t1134 517.045
R8457 VSS.t1497 VSS.t2085 517.045
R8458 VSS.t4020 VSS.t2528 517.045
R8459 VSS.t2000 VSS.t2486 517.045
R8460 VSS.t2967 VSS.t3173 517.045
R8461 VSS.t3274 VSS.t3967 517.045
R8462 VSS.t2071 VSS.t4227 517.045
R8463 VSS.t3939 VSS.t3217 517.045
R8464 VSS.t2408 VSS.t2506 517.045
R8465 VSS.t3016 VSS.t1189 517.045
R8466 VSS.t3478 VSS.t2618 517.045
R8467 VSS.t3807 VSS.t2116 517.045
R8468 VSS.t2779 VSS.t2847 517.045
R8469 VSS.t4237 VSS.t2264 517.045
R8470 VSS.t4233 VSS.t2357 517.045
R8471 VSS.t153 VSS.t1302 517.045
R8472 VSS.t1302 VSS.t157 517.045
R8473 VSS.t157 VSS.t1330 517.045
R8474 VSS.t1330 VSS.t155 517.045
R8475 VSS.t155 VSS.t4319 517.045
R8476 VSS.t4319 VSS.t151 517.045
R8477 VSS.t3804 VSS.t711 517.045
R8478 VSS.t114 VSS.t3804 517.045
R8479 VSS.t3870 VSS.t1891 517.045
R8480 VSS.t1259 VSS.t1610 517.045
R8481 VSS.t1443 VSS.t2482 517.045
R8482 VSS.t4330 VSS.t2209 517.045
R8483 VSS.t1658 VSS.t2819 517.045
R8484 VSS.t3336 VSS.t2067 517.045
R8485 VSS.t3215 VSS.t3782 517.045
R8486 VSS.n1329 VSS.t2986 517.045
R8487 VSS.t2563 VSS.t2250 517.045
R8488 VSS.t1994 VSS.t4026 517.045
R8489 VSS.t4170 VSS.t879 517.045
R8490 VSS.t1390 VSS.t1208 517.045
R8491 VSS.t2225 VSS.t4357 517.045
R8492 VSS.t3819 VSS.t3257 517.045
R8493 VSS.t3612 VSS.t3120 517.045
R8494 VSS.t2458 VSS.t3912 517.045
R8495 VSS.t3647 VSS.t3547 517.045
R8496 VSS.t3997 VSS.t1664 517.045
R8497 VSS.t3920 VSS.t2740 517.045
R8498 VSS.t2565 VSS.t3395 517.045
R8499 VSS.t1564 VSS.t3951 517.045
R8500 VSS.t3957 VSS.t1194 517.045
R8501 VSS.t3995 VSS.t1962 517.045
R8502 VSS.t2734 VSS.t3605 517.045
R8503 VSS.t2141 VSS.t1224 517.045
R8504 VSS.t1612 VSS.t3164 517.045
R8505 VSS.t1162 VSS.t4065 517.045
R8506 VSS.t2978 VSS.t2213 517.045
R8507 VSS.t4130 VSS.t1240 517.045
R8508 VSS.t2237 VSS.t4071 517.045
R8509 VSS.t820 VSS.t335 517.045
R8510 VSS.t1181 VSS.t2312 517.045
R8511 VSS.t2412 VSS.t3480 517.045
R8512 VSS.t4324 VSS.t1632 517.045
R8513 VSS.t3610 VSS.t4055 517.045
R8514 VSS.t2460 VSS.t971 517.045
R8515 VSS.t2112 VSS.t3852 517.045
R8516 VSS.t2533 VSS.t4346 517.045
R8517 VSS.t3680 VSS.t2252 517.045
R8518 VSS.t14 VSS.t2815 517.045
R8519 VSS.t408 VSS.t14 517.045
R8520 VSS.t2639 VSS.t3187 517.045
R8521 VSS.n1430 VSS.t1768 517.045
R8522 VSS.t4210 VSS.t981 517.045
R8523 VSS.t4079 VSS.t3908 517.045
R8524 VSS.t1312 VSS.t1153 517.045
R8525 VSS.t3589 VSS.t2542 512.429
R8526 VSS.t3184 VSS.t1231 512.429
R8527 VSS.t865 VSS.t3901 512.429
R8528 VSS.t1561 VSS.t2921 507.812
R8529 VSS.t3042 VSS.t511 503.197
R8530 VSS.t1248 VSS.t2219 503.197
R8531 VSS.t1580 VSS.t842 503.197
R8532 VSS.t2002 VSS.t3446 503.197
R8533 VSS.t1205 VSS.t1198 503.197
R8534 VSS.t1079 VSS.t1592 503.197
R8535 VSS.t799 VSS.t806 503.197
R8536 VSS.t1721 VSS.t2959 498.58
R8537 VSS.t1727 VSS.t3175 498.58
R8538 VSS.t1731 VSS.t4273 498.58
R8539 VSS.t1719 VSS.t990 498.58
R8540 VSS.t4269 VSS.t1234 498.58
R8541 VSS.t2275 VSS.t1749 498.58
R8542 VSS.t3281 VSS.t2630 498.58
R8543 VSS.n1333 VSS.t4160 498.58
R8544 VSS.t3500 VSS.t2188 498.58
R8545 VSS.t1411 VSS.t1696 498.58
R8546 VSS.n622 VSS.t2872 498.58
R8547 VSS.t539 VSS.n2126 485.94
R8548 VSS.t1797 VSS.t3637 484.731
R8549 VSS.t845 VSS.t3053 484.731
R8550 VSS.t3543 VSS.t3556 484.731
R8551 VSS.t3977 VSS.t1996 481.481
R8552 VSS.t1471 VSS.t3406 480.115
R8553 VSS.t3558 VSS.t3828 480.115
R8554 VSS.t747 VSS.t1096 480.115
R8555 VSS.t749 VSS.t1092 480.115
R8556 VSS.t133 VSS.t1207 480.115
R8557 VSS.t3643 VSS.t2776 480.115
R8558 VSS.t2878 VSS.t3419 480.115
R8559 VSS.t2299 VSS.t3383 480.115
R8560 VSS.t1761 VSS.t1910 475.498
R8561 VSS.t2338 VSS.t2155 475.498
R8562 VSS.t1447 VSS.t2450 475.498
R8563 VSS.t2480 VSS.t2452 475.498
R8564 VSS.t4180 VSS.t3838 470.882
R8565 VSS.t1802 VSS.t3955 470.882
R8566 VSS.t1856 VSS.t1299 470.882
R8567 VSS.t1160 VSS.t2692 466.264
R8568 VSS.t4116 VSS.t2660 466.264
R8569 VSS.t3545 VSS.t998 466.264
R8570 VSS.t2156 VSS.t2305 461.649
R8571 VSS.t319 VSS.t2617 461.649
R8572 VSS.t1535 VSS.t3138 461.649
R8573 VSS.t1688 VSS.t962 461.649
R8574 VSS.t2302 VSS.t1157 461.649
R8575 VSS.t3594 VSS.t2589 461.649
R8576 VSS.t2674 VSS.t3736 457.031
R8577 VSS.t2150 VSS.t1017 457.031
R8578 VSS.t1166 VSS.t303 457.031
R8579 VSS.t2950 VSS.t2668 457.031
R8580 VSS.t1904 VSS.t547 457.031
R8581 VSS.t2818 VSS.t3162 457.031
R8582 VSS.t2195 VSS.t1488 457.031
R8583 VSS.t2241 VSS.t797 457.031
R8584 VSS.t434 VSS.t4037 457.031
R8585 VSS.t3527 VSS.t3106 457.031
R8586 VSS.t2026 VSS.t2048 457.031
R8587 VSS.t1938 VSS.t3474 452.416
R8588 VSS.t3948 VSS.t4110 452.416
R8589 VSS.t1060 VSS.t899 447.798
R8590 VSS.t2567 VSS.t903 447.798
R8591 VSS.t3415 VSS.t3051 447.798
R8592 VSS.t3772 VSS.t3514 447.798
R8593 VSS.t1956 VSS.t674 443.183
R8594 VSS.t983 VSS.t1100 443.183
R8595 VSS.t2477 VSS.t1385 443.183
R8596 VSS.t634 VSS.n58 441.098
R8597 VSS.t97 VSS.n59 441.098
R8598 VSS.t1346 VSS.n60 441.098
R8599 VSS.t1822 VSS.n61 441.098
R8600 VSS.t248 VSS.n62 441.098
R8601 VSS.t587 VSS.n64 441.098
R8602 VSS.t719 VSS.n63 441.098
R8603 VSS.t741 VSS.n31 441.098
R8604 VSS.t1828 VSS.n32 441.098
R8605 VSS.t103 VSS.n33 441.098
R8606 VSS.t640 VSS.n34 441.098
R8607 VSS.t1352 VSS.n35 441.098
R8608 VSS.t254 VSS.n36 441.098
R8609 VSS.t575 VSS.n37 441.098
R8610 VSS.t3124 VSS.t3777 438.565
R8611 VSS.t2314 VSS.t1062 438.565
R8612 VSS.t4108 VSS.t1257 438.565
R8613 VSS.t2806 VSS.t34 438.565
R8614 VSS.n2456 VSS.t229 433.164
R8615 VSS.t2363 VSS.t2560 429.332
R8616 VSS.t3194 VSS.t773 429.332
R8617 VSS.t3278 VSS.t1487 429.332
R8618 VSS.t2178 VSS.t781 429.332
R8619 VSS.t3532 VSS.t4036 429.332
R8620 VSS.t183 VSS.t3300 424.716
R8621 VSS.t1168 VSS.t1309 424.716
R8622 VSS.t1220 VSS.t3865 424.716
R8623 VSS.t2046 VSS.t1072 424.716
R8624 VSS.t2990 VSS.t3352 424.716
R8625 VSS.t3742 VSS.t3438 424.716
R8626 VSS.t2520 VSS.t3542 420.099
R8627 VSS.t3760 VSS.t4049 420.099
R8628 VSS.t4040 VSS.t2352 420.099
R8629 VSS.t3385 VSS.t2924 420.099
R8630 VSS.t1509 VSS.t2522 420.099
R8631 VSS.t1041 VSS.t2270 415.483
R8632 VSS.t3607 VSS.n788 410.866
R8633 VSS.t1062 VSS.t1310 410.866
R8634 VSS.t4290 VSS.t2843 410.866
R8635 VSS.t2416 VSS.t1109 410.866
R8636 VSS.t3946 VSS.t983 406.25
R8637 VSS.t3442 VSS.t1709 401.635
R8638 VSS.t3795 VSS.t3862 401.635
R8639 VSS.t2537 VSS.t1569 397.017
R8640 VSS.t2602 VSS.t2220 397.017
R8641 VSS.t1629 VSS.t2114 397.017
R8642 VSS.t4110 VSS.t3676 397.017
R8643 VSS.t3082 VSS.t2674 392.401
R8644 VSS.t3684 VSS.t1570 392.401
R8645 VSS.t3897 VSS.t2150 392.401
R8646 VSS.t8 VSS.t817 392.401
R8647 VSS.t2029 VSS.t3898 392.401
R8648 VSS.t2643 VSS.t482 387.784
R8649 VSS.t4253 VSS.n856 387.784
R8650 VSS.t3943 VSS.t505 387.784
R8651 VSS.t1077 VSS.t767 383.168
R8652 VSS.t817 VSS.t1413 383.168
R8653 VSS.t3158 VSS.t2823 383.168
R8654 VSS.t3110 VSS.t3702 383.168
R8655 VSS.t1569 VSS.t2538 378.551
R8656 VSS.t2221 VSS.t2602 378.551
R8657 VSS.t2114 VSS.t1630 378.551
R8658 VSS.t3676 VSS.t4112 378.551
R8659 VSS.t1269 VSS.t521 373.935
R8660 VSS.t836 VSS.t1799 373.935
R8661 VSS.t1934 VSS.t1402 373.935
R8662 VSS.t40 VSS.t2708 373.935
R8663 VSS.t327 VSS.t787 369.318
R8664 VSS.t691 VSS.t3200 369.318
R8665 VSS.t526 VSS.t2169 369.318
R8666 VSS.t1850 VSS.t2106 369.318
R8667 VSS.t1604 VSS.t2688 369.318
R8668 VSS.t3575 VSS.t2217 369.318
R8669 VSS.t3724 VSS.t2682 369.318
R8670 VSS.t234 VSS.t840 369.318
R8671 VSS.t3571 VSS.t3447 369.318
R8672 VSS.t2813 VSS.t2684 369.318
R8673 VSS.t50 VSS.t4032 369.318
R8674 VSS.t52 VSS.t2676 369.318
R8675 VSS.t1118 VSS.t749 369.318
R8676 VSS.t3055 VSS.t133 369.318
R8677 VSS.t913 VSS.t1803 369.318
R8678 VSS.t911 VSS.t394 369.318
R8679 VSS.t800 VSS.t3373 369.318
R8680 VSS.t832 VSS.t392 369.318
R8681 VSS.t1670 VSS.t3436 369.318
R8682 VSS.t1674 VSS.t402 369.318
R8683 VSS.t916 VSS.t661 369.318
R8684 VSS.t400 VSS.t475 369.318
R8685 VSS.t4202 VSS.t4198 369.318
R8686 VSS.t803 VSS.t4200 369.318
R8687 VSS.t466 VSS.t3107 369.318
R8688 VSS.t2124 VSS.t4208 369.318
R8689 VSS.t3475 VSS.t1574 369.318
R8690 VSS.t3754 VSS.t826 364.786
R8691 VSS.t1982 VSS.t3361 364.702
R8692 VSS.t3053 VSS.t3316 364.702
R8693 VSS.n436 VSS.t4315 364.702
R8694 VSS.t3318 VSS.t3543 364.702
R8695 VSS.n2332 VSS.t4083 364.486
R8696 VSS.n527 VSS.t1795 360.587
R8697 VSS.t3927 VSS.t3320 355.469
R8698 VSS.t1954 VSS.t4147 355.469
R8699 VSS.t143 VSS.t4192 355.469
R8700 VSS.t2044 VSS.t4247 355.469
R8701 VSS.t1073 VSS.t4156 355.469
R8702 VSS.t694 VSS.t527 350.853
R8703 VSS.t3560 VSS.t1906 350.853
R8704 VSS.t1309 VSS.t1955 350.853
R8705 VSS.t1860 VSS.t295 350.853
R8706 VSS.t289 VSS.t1331 350.853
R8707 VSS.t1340 VSS.t2046 350.853
R8708 VSS.t869 VSS.t881 350.853
R8709 VSS.t859 VSS.t875 350.853
R8710 VSS.t861 VSS.t883 350.853
R8711 VSS.t2801 VSS.t650 350.853
R8712 VSS.t7 VSS.t3066 350.853
R8713 VSS.t513 VSS.t775 350.853
R8714 VSS.n2457 VSS.n2456 346.322
R8715 VSS.t2742 VSS.n980 346.236
R8716 VSS.t2664 VSS.t2532 346.236
R8717 VSS.t2268 VSS.t1969 343.279
R8718 VSS.n2455 VSS.n58 338.762
R8719 VSS.n2453 VSS.n59 338.762
R8720 VSS.n2451 VSS.n60 338.762
R8721 VSS.n2449 VSS.n61 338.762
R8722 VSS.n2447 VSS.n62 338.762
R8723 VSS.n2443 VSS.n64 338.762
R8724 VSS.n2445 VSS.n63 338.762
R8725 VSS.n2493 VSS.n31 338.762
R8726 VSS.n2493 VSS.n32 338.762
R8727 VSS.n2493 VSS.n33 338.762
R8728 VSS.n2493 VSS.n34 338.762
R8729 VSS.n2493 VSS.n35 338.762
R8730 VSS.n2493 VSS.n36 338.762
R8731 VSS.n2493 VSS.n37 338.762
R8732 VSS.t1231 VSS.t3295 337.003
R8733 VSS.t3779 VSS.t3124 337.003
R8734 VSS.t3944 VSS.t865 337.003
R8735 VSS.t34 VSS.t2805 337.003
R8736 VSS.t674 VSS.t1958 332.387
R8737 VSS.t3239 VSS.t1519 332.387
R8738 VSS.t9 VSS.t3670 332.387
R8739 VSS.t1149 VSS.t1897 332.387
R8740 VSS.t3868 VSS.t2077 332.387
R8741 VSS.t4075 VSS.t2073 332.387
R8742 VSS.t2722 VSS.t920 332.387
R8743 VSS.t959 VSS.t519 327.771
R8744 VSS.t3540 VSS.t1618 327.771
R8745 VSS.n2439 VSS.n2438 327.598
R8746 VSS.n2434 VSS.n2433 323.603
R8747 VSS.t1202 VSS.t398 323.154
R8748 VSS.t360 VSS.t1961 323.154
R8749 VSS.t919 VSS.t2195 318.538
R8750 VSS.t1466 VSS.t434 318.538
R8751 VSS.t3106 VSS.t3529 318.538
R8752 VSS.t2048 VSS.t2027 318.538
R8753 VSS.t3006 VSS.t2748 318.538
R8754 VSS.t1765 VSS.t2307 313.921
R8755 VSS.t1513 VSS.t3809 313.921
R8756 VSS.t2109 VSS.t3811 313.921
R8757 VSS.t3387 VSS.t3813 313.921
R8758 VSS.t1606 VSS.t4281 313.921
R8759 VSS.t1753 VSS.t2316 313.921
R8760 VSS.t509 VSS.t319 313.921
R8761 VSS.t2262 VSS.t1138 313.921
R8762 VSS.t3866 VSS.t432 313.921
R8763 VSS.t4030 VSS.t428 313.921
R8764 VSS.t2996 VSS.t46 313.921
R8765 VSS.t3152 VSS.t3574 313.921
R8766 VSS.t3578 VSS.t2590 313.921
R8767 VSS.t871 VSS.t3774 313.921
R8768 VSS.t3351 VSS.t607 313.921
R8769 VSS.t1805 VSS.t907 313.921
R8770 VSS.t1066 VSS.t905 313.921
R8771 VSS.t1865 VSS.t4206 313.921
R8772 VSS.t285 VSS.t3034 313.921
R8773 VSS.t3439 VSS.t1672 313.921
R8774 VSS.t3434 VSS.t1676 313.921
R8775 VSS.t3784 VSS.t1682 313.921
R8776 VSS.t1008 VSS.t177 313.921
R8777 VSS.t3299 VSS.t181 313.921
R8778 VSS.t4012 VSS.t3653 313.921
R8779 VSS.t821 VSS.t1688 313.921
R8780 VSS.t962 VSS.t2302 313.921
R8781 VSS.t3109 VSS.t3603 313.921
R8782 VSS.t4218 VSS.t930 313.921
R8783 VSS.t2692 VSS.t1159 309.305
R8784 VSS.t1445 VSS.t480 309.305
R8785 VSS.t3839 VSS.t4180 304.688
R8786 VSS.t26 VSS.t2087 304.688
R8787 VSS.t3734 VSS.t3127 304.688
R8788 VSS.n82 VSS.t1733 303.738
R8789 VSS.t761 VSS.t1083 303.156
R8790 VSS.t3849 VSS.t2338 300.072
R8791 VSS.t2998 VSS.t1334 300.072
R8792 VSS.t484 VSS.t2472 300.072
R8793 VSS.t1407 VSS.t3512 300.072
R8794 VSS.t1228 VSS.t4259 300.072
R8795 VSS.t1902 VSS.t2023 295.455
R8796 VSS.t3490 VSS.t1970 295.455
R8797 VSS.t3492 VSS.t918 295.455
R8798 VSS.t643 VSS.t1636 295.455
R8799 VSS.t4313 VSS.t3688 295.455
R8800 VSS.t937 VSS.n372 293.928
R8801 VSS.t3635 VSS.t1797 290.839
R8802 VSS.t823 VSS.t17 290.839
R8803 VSS.t1039 VSS.t504 286.223
R8804 VSS.t626 VSS.t613 282.303
R8805 VSS.t613 VSS.t632 282.303
R8806 VSS.t632 VSS.t622 282.303
R8807 VSS.t622 VSS.t641 282.303
R8808 VSS.t641 VSS.t620 282.303
R8809 VSS.t620 VSS.t636 282.303
R8810 VSS.t636 VSS.t628 282.303
R8811 VSS.t628 VSS.t615 282.303
R8812 VSS.t615 VSS.t634 282.303
R8813 VSS.t89 VSS.t76 282.303
R8814 VSS.t76 VSS.t95 282.303
R8815 VSS.t95 VSS.t85 282.303
R8816 VSS.t85 VSS.t74 282.303
R8817 VSS.t74 VSS.t83 282.303
R8818 VSS.t83 VSS.t99 282.303
R8819 VSS.t99 VSS.t91 282.303
R8820 VSS.t91 VSS.t78 282.303
R8821 VSS.t78 VSS.t97 282.303
R8822 VSS.t1368 VSS.t1355 282.303
R8823 VSS.t1355 VSS.t1344 282.303
R8824 VSS.t1344 VSS.t1364 282.303
R8825 VSS.t1364 VSS.t1353 282.303
R8826 VSS.t1353 VSS.t1362 282.303
R8827 VSS.t1362 VSS.t1348 282.303
R8828 VSS.t1348 VSS.t1370 282.303
R8829 VSS.t1370 VSS.t1357 282.303
R8830 VSS.t1357 VSS.t1346 282.303
R8831 VSS.t1844 VSS.t1831 282.303
R8832 VSS.t1831 VSS.t1820 282.303
R8833 VSS.t1820 VSS.t1840 282.303
R8834 VSS.t1840 VSS.t1829 282.303
R8835 VSS.t1829 VSS.t1838 282.303
R8836 VSS.t1838 VSS.t1824 282.303
R8837 VSS.t1824 VSS.t1846 282.303
R8838 VSS.t1846 VSS.t1833 282.303
R8839 VSS.t1833 VSS.t1822 282.303
R8840 VSS.t240 VSS.t257 282.303
R8841 VSS.t257 VSS.t246 282.303
R8842 VSS.t246 VSS.t266 282.303
R8843 VSS.t266 VSS.t255 282.303
R8844 VSS.t255 VSS.t264 282.303
R8845 VSS.t264 VSS.t250 282.303
R8846 VSS.t250 VSS.t242 282.303
R8847 VSS.t242 VSS.t259 282.303
R8848 VSS.t259 VSS.t248 282.303
R8849 VSS.t573 VSS.t601 282.303
R8850 VSS.t601 VSS.t567 282.303
R8851 VSS.t567 VSS.t585 282.303
R8852 VSS.t585 VSS.t597 282.303
R8853 VSS.t597 VSS.t569 282.303
R8854 VSS.t569 VSS.t591 282.303
R8855 VSS.t591 VSS.t603 282.303
R8856 VSS.t603 VSS.t577 282.303
R8857 VSS.t577 VSS.t587 282.303
R8858 VSS.t739 VSS.t729 282.303
R8859 VSS.t729 VSS.t734 282.303
R8860 VSS.t734 VSS.t717 282.303
R8861 VSS.t717 VSS.t726 282.303
R8862 VSS.t726 VSS.t736 282.303
R8863 VSS.t736 VSS.t722 282.303
R8864 VSS.t722 VSS.t731 282.303
R8865 VSS.t731 VSS.t742 282.303
R8866 VSS.t742 VSS.t719 282.303
R8867 VSS.t728 VSS.t745 282.303
R8868 VSS.t745 VSS.t724 282.303
R8869 VSS.t724 VSS.t733 282.303
R8870 VSS.t733 VSS.t744 282.303
R8871 VSS.t744 VSS.t721 282.303
R8872 VSS.t721 VSS.t738 282.303
R8873 VSS.t738 VSS.t746 282.303
R8874 VSS.t746 VSS.t725 282.303
R8875 VSS.t725 VSS.t741 282.303
R8876 VSS.t1835 VSS.t1837 282.303
R8877 VSS.t1837 VSS.t1827 282.303
R8878 VSS.t1827 VSS.t1848 282.303
R8879 VSS.t1848 VSS.t1836 282.303
R8880 VSS.t1836 VSS.t1826 282.303
R8881 VSS.t1826 VSS.t1843 282.303
R8882 VSS.t1843 VSS.t1849 282.303
R8883 VSS.t1849 VSS.t1842 282.303
R8884 VSS.t1842 VSS.t1828 282.303
R8885 VSS.t80 VSS.t82 282.303
R8886 VSS.t82 VSS.t102 282.303
R8887 VSS.t102 VSS.t93 282.303
R8888 VSS.t93 VSS.t81 282.303
R8889 VSS.t81 VSS.t101 282.303
R8890 VSS.t101 VSS.t88 282.303
R8891 VSS.t88 VSS.t94 282.303
R8892 VSS.t94 VSS.t87 282.303
R8893 VSS.t87 VSS.t103 282.303
R8894 VSS.t617 VSS.t619 282.303
R8895 VSS.t619 VSS.t639 282.303
R8896 VSS.t639 VSS.t630 282.303
R8897 VSS.t630 VSS.t618 282.303
R8898 VSS.t618 VSS.t638 282.303
R8899 VSS.t638 VSS.t625 282.303
R8900 VSS.t625 VSS.t631 282.303
R8901 VSS.t631 VSS.t624 282.303
R8902 VSS.t624 VSS.t640 282.303
R8903 VSS.t1359 VSS.t1361 282.303
R8904 VSS.t1361 VSS.t1351 282.303
R8905 VSS.t1351 VSS.t1372 282.303
R8906 VSS.t1372 VSS.t1360 282.303
R8907 VSS.t1360 VSS.t1350 282.303
R8908 VSS.t1350 VSS.t1367 282.303
R8909 VSS.t1367 VSS.t1373 282.303
R8910 VSS.t1373 VSS.t1366 282.303
R8911 VSS.t1366 VSS.t1352 282.303
R8912 VSS.t261 VSS.t263 282.303
R8913 VSS.t263 VSS.t253 282.303
R8914 VSS.t253 VSS.t244 282.303
R8915 VSS.t244 VSS.t262 282.303
R8916 VSS.t262 VSS.t252 282.303
R8917 VSS.t252 VSS.t239 282.303
R8918 VSS.t239 VSS.t245 282.303
R8919 VSS.t245 VSS.t268 282.303
R8920 VSS.t268 VSS.t254 282.303
R8921 VSS.t599 VSS.t581 282.303
R8922 VSS.t581 VSS.t593 282.303
R8923 VSS.t593 VSS.t605 282.303
R8924 VSS.t605 VSS.t579 282.303
R8925 VSS.t579 VSS.t589 282.303
R8926 VSS.t589 VSS.t571 282.303
R8927 VSS.t571 VSS.t583 282.303
R8928 VSS.t583 VSS.t595 282.303
R8929 VSS.t595 VSS.t575 282.303
R8930 VSS.t2628 VSS.t3281 276.99
R8931 VSS.t751 VSS.t1094 276.99
R8932 VSS.t2186 VSS.t3500 276.99
R8933 VSS.t2219 VSS.t1249 272.373
R8934 VSS.t502 VSS.t2161 272.373
R8935 VSS.t3446 VSS.t2003 272.373
R8936 VSS.t3822 VSS.t1087 267.757
R8937 VSS.t857 VSS.t856 267.49
R8938 VSS.t1997 VSS.t3977 267.49
R8939 VSS.t2500 VSS.t2451 267.49
R8940 VSS.t3776 VSS.t2088 264.687
R8941 VSS.t2542 VSS.t3590 263.139
R8942 VSS.t2318 VSS.t189 263.139
R8943 VSS.t1229 VSS.t3184 263.139
R8944 VSS.t1187 VSS.t2612 263.139
R8945 VSS.t3657 VSS.t2916 258.524
R8946 VSS.t2021 VSS.t3261 258.524
R8947 VSS.t2947 VSS.t1014 258.524
R8948 VSS.t1025 VSS.t3001 258.524
R8949 VSS.t151 VSS.t2826 258.524
R8950 VSS.t139 VSS.t3473 258.524
R8951 VSS.t137 VSS.t3472 258.524
R8952 VSS.t1208 VSS.t1389 258.524
R8953 VSS.t2426 VSS.t2383 258.236
R8954 VSS.t235 VSS.t937 256.137
R8955 VSS.t1431 VSS.n379 256.137
R8956 VSS.t1576 VSS.t1518 253.906
R8957 VSS.t1091 VSS.t3597 253.906
R8958 VSS.t3168 VSS.t2922 249.291
R8959 VSS.t4083 VSS.t2943 245.161
R8960 VSS.t3667 VSS.t1877 244.673
R8961 VSS.t1862 VSS.t3516 244.673
R8962 VSS.t1064 VSS.t3780 242.992
R8963 VSS.t4229 VSS.t1064 242.992
R8964 VSS.t3592 VSS.t4229 242.992
R8965 VSS.t2398 VSS.t3592 242.992
R8966 VSS.t3576 VSS.t2398 242.992
R8967 VSS.t4118 VSS.t3576 242.992
R8968 VSS.t4249 VSS.t4118 242.992
R8969 VSS.t3291 VSS.t1623 242.992
R8970 VSS.t1623 VSS.t2340 242.992
R8971 VSS.t2340 VSS.t2404 242.992
R8972 VSS.t2404 VSS.t4053 242.992
R8973 VSS.t4053 VSS.t3802 242.992
R8974 VSS.t3802 VSS.t2787 242.992
R8975 VSS.t2787 VSS.t2464 242.992
R8976 VSS.t3455 VSS.t3378 242.992
R8977 VSS.t3378 VSS.t3910 242.992
R8978 VSS.t3910 VSS.t4174 242.992
R8979 VSS.t4174 VSS.t3092 242.992
R8980 VSS.t3092 VSS.t1521 242.992
R8981 VSS.t1521 VSS.t2912 242.992
R8982 VSS.t2912 VSS.t1523 242.992
R8983 VSS.t2053 VSS.t3114 242.992
R8984 VSS.t3800 VSS.t2053 242.992
R8985 VSS.t1818 VSS.t3800 242.992
R8986 VSS.t2324 VSS.t1818 242.992
R8987 VSS.t2919 VSS.t2324 242.992
R8988 VSS.t2135 VSS.t2919 242.992
R8989 VSS.t3798 VSS.t2135 242.992
R8990 VSS.t2474 VSS.t2620 242.992
R8991 VSS.t4326 VSS.t2474 242.992
R8992 VSS.t3358 VSS.t4326 242.992
R8993 VSS.t1582 VSS.t3358 242.992
R8994 VSS.t1381 VSS.t1582 242.992
R8995 VSS.t2849 VSS.t1381 242.992
R8996 VSS.t4085 VSS.t2849 242.992
R8997 VSS.t2088 VSS.t3020 242.992
R8998 VSS.t3020 VSS.t4081 242.992
R8999 VSS.t4081 VSS.t3204 242.992
R9000 VSS.t3428 VSS.t126 240.058
R9001 VSS.t3732 VSS.t1621 240.058
R9002 VSS.t804 VSS.t2406 240.058
R9003 VSS.t949 VSS.t2143 239.341
R9004 VSS.t3375 VSS.t2171 235.44
R9005 VSS.t537 VSS.t1276 235.44
R9006 VSS.t1503 VSS.t2817 235.44
R9007 VSS.t3595 VSS.t3193 235.44
R9008 VSS.t1528 VSS.t3276 235.44
R9009 VSS.t4003 VSS.t2177 235.44
R9010 VSS.t1641 VSS.t3530 235.44
R9011 VSS.t2010 VSS.t1784 235.143
R9012 VSS.t450 VSS.t1690 235.143
R9013 VSS.t4102 VSS.t3990 235.143
R9014 VSS.t826 VSS.t769 235.143
R9015 VSS.t1280 VSS.t1948 230.825
R9016 VSS.t4182 VSS.t3830 230.825
R9017 VSS.t498 VSS.t838 226.208
R9018 VSS.t1859 VSS.t3686 226.208
R9019 VSS.t2732 VSS.t2206 226.208
R9020 VSS.t3063 VSS.t1449 226.208
R9021 VSS.n865 VSS.t1989 221.591
R9022 VSS.t21 VSS.t2606 221.591
R9023 VSS.t3169 VSS.t2860 221.591
R9024 VSS.t1733 VSS.t941 221.296
R9025 VSS.t2744 VSS.t2810 216.975
R9026 VSS.t420 VSS.t1578 216.975
R9027 VSS.t1875 VSS.t3549 216.975
R9028 VSS.t1531 VSS.t789 216.975
R9029 VSS.t3279 VSS.t1274 216.975
R9030 VSS.t1628 VSS.t352 216.975
R9031 VSS.t783 VSS.t3314 216.975
R9032 VSS.t3461 VSS.t3770 216.975
R9033 VSS.t2580 VSS.t1122 216.975
R9034 VSS.t1572 VSS.t3706 216.975
R9035 VSS.n2457 VSS.t216 212.53
R9036 VSS.t2627 VSS.t11 212.358
R9037 VSS.t647 VSS.t1105 212.358
R9038 VSS.t854 VSS.t657 212.358
R9039 VSS.n2492 VSS.t222 211.921
R9040 VSS.t2367 VSS.t1657 207.742
R9041 VSS.t2930 VSS.t2715 207.742
R9042 VSS.t851 VSS.t2982 207.742
R9043 VSS.t2280 VSS.t2498 207.742
R9044 VSS.n2421 VSS.t698 206.108
R9045 VSS.t3587 VSS.t4142 203.125
R9046 VSS.t4061 VSS.t3557 203.125
R9047 VSS.t688 VSS.t3026 203.125
R9048 VSS.t317 VSS.t1 203.125
R9049 VSS.t311 VSS.t2274 203.125
R9050 VSS.t309 VSS.t1625 203.125
R9051 VSS.t1263 VSS.t2649 203.125
R9052 VSS.t423 VSS.t4348 203.125
R9053 VSS.t1132 VSS.t540 203.125
R9054 VSS.t3756 VSS.t48 203.125
R9055 VSS.t426 VSS.t549 203.125
R9056 VSS.t163 VSS.t493 203.125
R9057 VSS.t161 VSS.t4194 203.125
R9058 VSS.t145 VSS.t812 203.125
R9059 VSS.t3328 VSS.t4114 203.125
R9060 VSS.t2266 VSS.t3858 203.125
R9061 VSS.t3330 VSS.t1328 203.125
R9062 VSS.t3045 VSS.t609 203.125
R9063 VSS.t611 VSS.t517 203.125
R9064 VSS.t500 VSS.t1854 203.125
R9065 VSS.t3008 VSS.t1684 203.125
R9066 VSS.t1678 VSS.t553 203.125
R9067 VSS.t173 VSS.t801 203.125
R9068 VSS.t963 VSS.t175 203.125
R9069 VSS.t792 VSS.t2517 203.125
R9070 VSS.t753 VSS.t1416 203.125
R9071 VSS.t1485 VSS.t328 203.125
R9072 VSS.t3310 VSS.t1147 203.125
R9073 VSS.n578 VSS.n577 202.722
R9074 VSS.t1793 VSS.n526 197.351
R9075 VSS.t1454 VSS.t333 193.893
R9076 VSS.t4190 VSS.t3342 193.893
R9077 VSS.t2 VSS.t3130 193.678
R9078 VSS.t3864 VSS.n2125 189.276
R9079 VSS.t4311 VSS.t2223 184.66
R9080 VSS.t4307 VSS.t2387 184.66
R9081 VSS.t1056 VSS.t3655 184.66
R9082 VSS.t1048 VSS.t3786 184.66
R9083 VSS.t1044 VSS.t1694 184.66
R9084 VSS.t1052 VSS.t3057 184.66
R9085 VSS.t825 VSS.t2137 184.66
R9086 VSS.t2079 VSS.t1272 184.66
R9087 VSS.t1600 VSS.t2055 184.66
R9088 VSS.t3453 VSS.t532 184.66
R9089 VSS.t2065 VSS.t795 184.66
R9090 VSS.t3208 VSS.t1899 184.66
R9091 VSS.t645 VSS.n708 184.66
R9092 VSS.t1314 VSS.t2868 184.66
R9093 VSS.t32 VSS.t2096 184.66
R9094 VSS.t3878 VSS.t1660 184.66
R9095 VSS.t2344 VSS.t2738 184.66
R9096 VSS.n2233 VSS.n2232 184.413
R9097 VSS.t3780 VSS.n2233 182.244
R9098 VSS.n2234 VSS.t4249 182.244
R9099 VSS.n2234 VSS.t3291 182.244
R9100 VSS.t2464 VSS.n90 182.244
R9101 VSS.n90 VSS.t3455 182.244
R9102 VSS.n2330 VSS.t1523 182.244
R9103 VSS.t3114 VSS.n2330 182.244
R9104 VSS.n2331 VSS.t3798 182.244
R9105 VSS.t2620 VSS.n2331 182.244
R9106 VSS.n2332 VSS.t4085 182.244
R9107 VSS.t3204 VSS.n82 182.244
R9108 VSS.t2290 VSS.t1322 180.043
R9109 VSS.t867 VSS.t1858 180.043
R9110 VSS.t901 VSS.t3609 180.043
R9111 VSS.t810 VSS.t1879 180.043
R9112 VSS.t1541 VSS.t852 180.043
R9113 VSS.n2217 VSS.n372 178.457
R9114 VSS.n486 VSS.t1546 178.457
R9115 VSS.t3523 VSS.n504 178.457
R9116 VSS.t648 VSS.t858 178.327
R9117 VSS.t855 VSS.t1107 176.903
R9118 VSS.n505 VSS.t3482 174.257
R9119 VSS.t2144 VSS.t3754 173.208
R9120 VSS.t2365 VSS.t2562 170.81
R9121 VSS.t3614 VSS.t2396 170.81
R9122 VSS.t171 VSS.t3831 170.81
R9123 VSS.t3170 VSS.t4162 170.81
R9124 VSS.t1006 VSS.t3346 170.81
R9125 VSS.t545 VSS.t3401 170.81
R9126 VSS.t1999 VSS.t3399 170.81
R9127 VSS.t477 VSS.t2377 166.194
R9128 VSS.t3572 VSS.t3999 166.194
R9129 VSS.t3360 VSS.t2034 166.194
R9130 VSS.n984 VSS.t2108 166.194
R9131 VSS.t3926 VSS.t4137 166.194
R9132 VSS.t299 VSS.t686 166.194
R9133 VSS.t297 VSS.t4063 166.194
R9134 VSS.t507 VSS.t1483 166.194
R9135 VSS.t281 VSS.t165 166.194
R9136 VSS.t1332 VSS.t169 166.194
R9137 VSS.t358 VSS.t3918 166.194
R9138 VSS.t2133 VSS.t3580 166.194
R9139 VSS.t3642 VSS.n644 166.194
R9140 VSS.t1119 VSS.t2125 166.194
R9141 VSS.t4092 VSS.t813 166.194
R9142 VSS.t15 VSS.t4104 166.194
R9143 VSS.t2822 VSS.t13 166.194
R9144 VSS.t3961 VSS.t816 166.194
R9145 VSS.t4295 VSS.t2581 166.194
R9146 VSS.t1155 VSS.t2862 166.194
R9147 VSS.n2493 VSS.n2492 162.755
R9148 VSS.t3758 VSS.t4048 161.577
R9149 VSS.t1101 VSS.t3030 161.577
R9150 VSS.t3947 VSS.t3599 161.577
R9151 VSS.n486 VSS.t710 159.036
R9152 VSS.n541 VSS.t3845 157.462
R9153 VSS.n379 VSS.t2573 155.363
R9154 VSS.n504 VSS.t1741 155.363
R9155 VSS.n505 VSS.t1173 155.363
R9156 VSS.n526 VSS.t2795 155.363
R9157 VSS.n527 VSS.t2420 155.363
R9158 VSS.t4136 VSS.t5 152.345
R9159 VSS.t3117 VSS.t1376 152.345
R9160 VSS.t2414 VSS.t3696 152.345
R9161 VSS.t2050 VSS.t44 152.345
R9162 VSS.t2272 VSS.t321 147.727
R9163 VSS.t2686 VSS.t307 147.727
R9164 VSS.t516 VSS.t1068 147.727
R9165 VSS.t3716 VSS.t915 147.119
R9166 VSS.t2943 VSS.t3466 141.022
R9167 VSS.t3482 VSS.t4102 140.666
R9168 VSS.t3466 VSS.t3776 138.852
R9169 VSS.t755 VSS.t1121 138.494
R9170 VSS.t1546 VSS.t2010 136.466
R9171 VSS.t1690 VSS.t3523 136.466
R9172 VSS.t2383 VSS.t3845 136.466
R9173 VSS.t208 VSS.t225 136.019
R9174 VSS.t225 VSS.t214 136.019
R9175 VSS.t214 VSS.t204 136.019
R9176 VSS.t204 VSS.t223 136.019
R9177 VSS.t223 VSS.t202 136.019
R9178 VSS.t202 VSS.t218 136.019
R9179 VSS.t218 VSS.t210 136.019
R9180 VSS.t210 VSS.t227 136.019
R9181 VSS.t227 VSS.t216 136.019
R9182 VSS.t229 VSS.t231 135.63
R9183 VSS.t231 VSS.t221 135.63
R9184 VSS.t221 VSS.t212 135.63
R9185 VSS.t212 VSS.t230 135.63
R9186 VSS.t230 VSS.t220 135.63
R9187 VSS.t220 VSS.t207 135.63
R9188 VSS.t207 VSS.t213 135.63
R9189 VSS.t213 VSS.t206 135.63
R9190 VSS.t206 VSS.t222 135.63
R9191 VSS.t769 VSS.t1793 134.368
R9192 VSS.t3494 VSS.t1971 133.879
R9193 VSS.t3496 VSS.t2980 133.879
R9194 VSS.t765 VSS.t4263 133.879
R9195 VSS.t849 VSS.t2874 133.879
R9196 VSS.t2031 VSS.t1792 133.879
R9197 VSS.n2431 VSS.n2430 133.835
R9198 VSS.t1255 VSS.n764 129.262
R9199 VSS.t2090 VSS.t491 129.262
R9200 VSS.t2254 VSS.t808 129.262
R9201 VSS.n577 VSS.t374 126.612
R9202 VSS.t706 VSS.t24 124.829
R9203 VSS.t704 VSS.t25 124.829
R9204 VSS.t4245 VSS.t2199 124.645
R9205 VSS.t4115 VSS.t987 124.645
R9206 VSS.n648 VSS.t3322 124.645
R9207 VSS.t1126 VSS.t1594 124.645
R9208 VSS.t1113 VSS.t1596 124.645
R9209 VSS.t2821 VSS.t1929 124.645
R9210 VSS.t941 VSS.t939 121.496
R9211 VSS.t939 VSS.t945 121.496
R9212 VSS.t945 VSS.t943 121.496
R9213 VSS.t943 VSS.t669 121.496
R9214 VSS.t669 VSS.t667 121.496
R9215 VSS.t667 VSS.t696 121.496
R9216 VSS.t696 VSS.t715 121.496
R9217 VSS.t715 VSS.t700 121.496
R9218 VSS.t700 VSS.t671 121.496
R9219 VSS.t671 VSS.t713 121.496
R9220 VSS.t713 VSS.t698 121.496
R9221 VSS.t237 VSS.t235 117.572
R9222 VSS.t275 VSS.t237 117.572
R9223 VSS.t279 VSS.t275 117.572
R9224 VSS.t271 VSS.t279 117.572
R9225 VSS.t273 VSS.t271 117.572
R9226 VSS.t277 VSS.t273 117.572
R9227 VSS.t269 VSS.t277 117.572
R9228 VSS.t2571 VSS.t269 117.572
R9229 VSS.t2577 VSS.t2571 117.572
R9230 VSS.t2575 VSS.t2577 117.572
R9231 VSS.t2573 VSS.t2575 117.572
R9232 VSS.t1437 VSS.t1431 117.572
R9233 VSS.t1429 VSS.t1437 117.572
R9234 VSS.t1441 VSS.t1429 117.572
R9235 VSS.t1435 VSS.t1441 117.572
R9236 VSS.t1427 VSS.t1435 117.572
R9237 VSS.t1433 VSS.t1427 117.572
R9238 VSS.t1439 VSS.t1433 117.572
R9239 VSS.t3134 VSS.t1439 117.572
R9240 VSS.t3132 VSS.t3134 117.572
R9241 VSS.t3136 VSS.t3132 117.572
R9242 VSS.t3130 VSS.t3136 117.572
R9243 VSS.t1784 VSS.t1790 117.572
R9244 VSS.t1790 VSS.t1780 117.572
R9245 VSS.t1780 VSS.t1776 117.572
R9246 VSS.t1776 VSS.t1788 117.572
R9247 VSS.t1788 VSS.t1782 117.572
R9248 VSS.t1782 VSS.t1786 117.572
R9249 VSS.t1786 VSS.t1778 117.572
R9250 VSS.t1778 VSS.t1737 117.572
R9251 VSS.t1737 VSS.t1735 117.572
R9252 VSS.t1735 VSS.t1739 117.572
R9253 VSS.t1739 VSS.t1741 117.572
R9254 VSS.t442 VSS.t450 117.572
R9255 VSS.t448 VSS.t442 117.572
R9256 VSS.t436 VSS.t448 117.572
R9257 VSS.t440 VSS.t436 117.572
R9258 VSS.t446 VSS.t440 117.572
R9259 VSS.t438 VSS.t446 117.572
R9260 VSS.t444 VSS.t438 117.572
R9261 VSS.t1175 VSS.t444 117.572
R9262 VSS.t1171 VSS.t1175 117.572
R9263 VSS.t1169 VSS.t1171 117.572
R9264 VSS.t1173 VSS.t1169 117.572
R9265 VSS.t3990 VSS.t3982 117.572
R9266 VSS.t3982 VSS.t3988 117.572
R9267 VSS.t3988 VSS.t3992 117.572
R9268 VSS.t3992 VSS.t3980 117.572
R9269 VSS.t3980 VSS.t3986 117.572
R9270 VSS.t3986 VSS.t3978 117.572
R9271 VSS.t3978 VSS.t3984 117.572
R9272 VSS.t3984 VSS.t2789 117.572
R9273 VSS.t2789 VSS.t2793 117.572
R9274 VSS.t2793 VSS.t2791 117.572
R9275 VSS.t2791 VSS.t2795 117.572
R9276 VSS.t1795 VSS.t950 117.572
R9277 VSS.t2420 VSS.t2440 117.572
R9278 VSS.t2440 VSS.t2442 117.572
R9279 VSS.t2442 VSS.t2438 117.572
R9280 VSS.t2438 VSS.t2436 117.572
R9281 VSS.t2436 VSS.t2424 117.572
R9282 VSS.t2424 VSS.t2432 117.572
R9283 VSS.t2432 VSS.t2434 117.572
R9284 VSS.t2434 VSS.t2428 117.572
R9285 VSS.t2428 VSS.t2430 117.572
R9286 VSS.t2430 VSS.t2422 117.572
R9287 VSS.t2422 VSS.t2426 117.572
R9288 VSS.t4038 VSS.n1994 115.412
R9289 VSS.n636 VSS.t1196 115.412
R9290 VSS.t1932 VSS.t1403 115.412
R9291 VSS.t3049 VSS.t2609 115.412
R9292 VSS.t28 VSS.t2841 115.412
R9293 VSS.t30 VSS.t2709 115.412
R9294 VSS.t4292 VSS.t3914 115.412
R9295 VSS.t338 VSS.n2549 111.499
R9296 VSS.t378 VSS.n48 106.936
R9297 VSS.t2599 VSS.t935 106.18
R9298 VSS.t2244 VSS.t3365 106.18
R9299 VSS.t926 VSS.t2342 106.18
R9300 VSS.n2422 VSS.n2421 105.225
R9301 VSS.n542 VSS.n541 101.826
R9302 VSS.t3836 VSS.t679 101.562
R9303 VSS.t1415 VSS.t3219 96.9465
R9304 VSS.t710 VSS.t2 96.5767
R9305 VSS.t1408 VSS.t3674 92.33
R9306 VSS.t1711 VSS.t3432 92.33
R9307 VSS.t0 VSS.t1747 92.33
R9308 VSS.t2582 VSS.t3720 92.33
R9309 VSS.n2519 VSS.n2516 89.2711
R9310 VSS.t2143 VSS.t2144 88.1788
R9311 VSS.t950 VSS.t949 88.1788
R9312 VSS.t933 VSS.t487 87.7136
R9313 VSS.t4361 VSS.t4073 87.7136
R9314 VSS.t2666 VSS.t2530 87.7136
R9315 VSS.t4221 VSS.t1383 87.7136
R9316 VSS.t3221 VSS.t1417 87.7136
R9317 VSS.t655 VSS.t785 87.7136
R9318 VSS.t396 VSS.t815 83.9154
R9319 VSS.n2526 VSS.n2514 83.8639
R9320 VSS.t3270 VSS.n905 83.0971
R9321 VSS.n2443 VSS.n2442 82.9471
R9322 VSS.n2445 VSS.n2444 82.9471
R9323 VSS.n2447 VSS.n2446 82.9471
R9324 VSS.n2449 VSS.n2448 82.9471
R9325 VSS.n2451 VSS.n2450 82.9471
R9326 VSS.n2453 VSS.n2452 82.9471
R9327 VSS.n2455 VSS.n2454 82.9471
R9328 VSS.t2092 VSS.n2523 82.6977
R9329 VSS.n2533 VSS.t3091 82.6977
R9330 VSS.n2548 VSS.t1400 82.4713
R9331 VSS.t4106 VSS.t3797 78.4806
R9332 VSS.t287 VSS.t2291 78.4806
R9333 VSS.t19 VSS.t1542 78.4806
R9334 VSS.t135 VSS.t16 73.8641
R9335 VSS.n2539 VSS.n2512 71.9895
R9336 VSS.t330 VSS.n2515 71.4594
R9337 VSS.t3212 VSS.t1620 69.2477
R9338 VSS.t2977 VSS.t1075 69.2477
R9339 VSS.t3069 VSS.n1451 69.2477
R9340 VSS.t846 VSS.t3430 69.2477
R9341 VSS.t3692 VSS.t3708 69.2477
R9342 VSS.t374 VSS.t376 68.4396
R9343 VSS.t376 VSS.t380 68.4396
R9344 VSS.t380 VSS.t382 68.4396
R9345 VSS.t382 VSS.t386 68.4396
R9346 VSS.t386 VSS.t390 68.4396
R9347 VSS.t390 VSS.t384 68.4396
R9348 VSS.t384 VSS.t388 68.4396
R9349 VSS.t388 VSS.t372 68.4396
R9350 VSS.t372 VSS.t378 68.4396
R9351 VSS.t1204 VSS.t362 64.6312
R9352 VSS.t331 VSS.t1452 64.6312
R9353 VSS.t368 VSS.t1959 64.6312
R9354 VSS.n2513 VSS.t897 60.4331
R9355 VSS.t3698 VSS.t2373 60.0147
R9356 VSS.t4316 VSS.t2129 60.0147
R9357 VSS.t2336 VSS.t2051 55.3982
R9358 VSS.t2519 VSS.t3815 55.3982
R9359 VSS.t3718 VSS.t676 55.3982
R9360 VSS.t3266 VSS.t430 55.3982
R9361 VSS.t1887 VSS.t3140 55.3982
R9362 VSS.t3079 VSS.t4215 55.3982
R9363 VSS.t3410 VSS.t909 55.3982
R9364 VSS.t2954 VSS.t1680 55.3982
R9365 VSS.t3301 VSS.t185 55.3982
R9366 VSS.t457 VSS.n2513 54.9199
R9367 VSS.t1082 VSS.t708 53.4984
R9368 VSS.t1655 VSS.t2371 50.7817
R9369 VSS.t3969 VSS.t1267 50.7817
R9370 VSS.t2904 VSS.t3823 50.7817
R9371 VSS.t2713 VSS.t1325 50.7817
R9372 VSS.t759 VSS.t18 46.1653
R9373 VSS.t1084 VSS.t757 45.3599
R9374 VSS.n2494 VSS.n2493 40.1356
R9375 VSS.t4289 VSS.t2641 36.9323
R9376 VSS.t2007 VSS.t3941 36.9323
R9377 VSS.t4098 VSS.t1553 36.9323
R9378 VSS.t1115 VSS.n715 36.9323
R9379 VSS.t4100 VSS.t649 36.9323
R9380 VSS.t64 VSS.n2494 35.1056
R9381 VSS.n2549 VSS.t1398 34.896
R9382 VSS.t486 VSS.t2611 32.3158
R9383 VSS.t2036 VSS.t2315 32.3158
R9384 VSS.t3183 VSS.t3151 32.3158
R9385 VSS.t1451 VSS.t4204 32.3158
R9386 VSS.t2094 VSS.n2515 31.5951
R9387 VSS.n2540 VSS.n2539 30.6409
R9388 VSS.n2524 VSS.n2514 28.7325
R9389 VSS.t2914 VSS.t1700 27.6994
R9390 VSS.t1320 VSS.t3882 27.6994
R9391 VSS.t1318 VSS.t2296 27.6994
R9392 VSS.n2540 VSS.t1400 26.506
R9393 VSS.t897 VSS.n2512 26.506
R9394 VSS.n2526 VSS.t457 26.506
R9395 VSS.n2524 VSS.t2092 26.506
R9396 VSS.n2523 VSS.t2094 26.506
R9397 VSS.n2519 VSS.t330 26.506
R9398 VSS.n2517 VSS.t3091 26.506
R9399 VSS.t2083 VSS.n2533 26.506
R9400 VSS.t1398 VSS.n2548 26.1983
R9401 VSS.t2624 VSS.t844 23.0829
R9402 VSS.t839 VSS.t2512 23.0829
R9403 VSS.t1816 VSS.t3377 23.0829
R9404 VSS.n915 VSS.t1811 18.4664
R9405 VSS.n921 VSS.t1568 18.4664
R9406 VSS.t3171 VSS.t692 18.4664
R9407 VSS.t1218 VSS.t4031 18.4664
R9408 VSS.t4168 VSS.t1511 18.4664
R9409 VSS.t4166 VSS.t3824 18.4664
R9410 VSS.t2992 VSS.t1806 18.4664
R9411 VSS.t3748 VSS.t3435 18.4664
R9412 VSS.t187 VSS.t1011 18.4664
R9413 VSS.n614 VSS.t3470 18.4664
R9414 VSS.t58 VSS.t344 15.6144
R9415 VSS.t70 VSS.t346 15.6144
R9416 VSS.t56 VSS.t342 15.6144
R9417 VSS.t68 VSS.t348 15.6144
R9418 VSS.t62 VSS.t350 15.6144
R9419 VSS.t54 VSS.t354 15.6144
R9420 VSS.t66 VSS.t356 15.6144
R9421 VSS.t60 VSS.t340 15.6144
R9422 VSS.t72 VSS.t336 15.6144
R9423 VSS.t1304 VSS.t1767 13.8499
R9424 VSS.t1216 VSS.t1058 13.8499
R9425 VSS.t1627 VSS.t2047 13.8499
R9426 VSS.t3585 VSS.t496 13.8499
R9427 VSS.t2994 VSS.t1936 13.8499
R9428 VSS.t3746 VSS.t3633 13.8499
R9429 VSS.t4265 VSS.t3369 13.8499
R9430 VSS.t819 VSS.t827 13.8499
R9431 VSS.t2588 VSS.t654 13.8499
R9432 VSS.n1012 VSS.t2545 11.0252
R9433 VSS.n1002 VSS.t3388 11.0252
R9434 VSS.n954 VSS.t1762 11.0252
R9435 VSS.n935 VSS.t1607 11.0252
R9436 VSS.n964 VSS.t1472 11.0252
R9437 VSS.n1847 VSS.t3027 11.0252
R9438 VSS.n1865 VSS.t1626 11.0252
R9439 VSS.n879 VSS.t2263 11.0252
R9440 VSS.n1899 VSS.t2931 11.0252
R9441 VSS.n813 VSS.t2997 11.0252
R9442 VSS.n1983 VSS.t1880 11.0252
R9443 VSS.n2006 VSS.t970 11.0252
R9444 VSS.n1975 VSS.t1303 11.0252
R9445 VSS.n731 VSS.t1585 11.0252
R9446 VSS.n703 VSS.t2861 11.0252
R9447 VSS.n667 VSS.t1067 11.0252
R9448 VSS.n2053 VSS.t22 11.0252
R9449 VSS.n1470 VSS.t3386 11.0252
R9450 VSS.n2156 VSS.t1855 11.0252
R9451 VSS.n571 VSS.t3785 11.0252
R9452 VSS.n2160 VSS.t4105 11.0252
R9453 VSS.n387 VSS.t3962 11.0252
R9454 VSS.n2180 VSS.t2518 11.0252
R9455 VSS.n451 VSS.t1697 11.0252
R9456 VSS.n595 VSS.t4043 11.0252
R9457 VSS.n586 VSS.t1637 11.0252
R9458 VSS.n2194 VSS.t2551 11.0252
R9459 VSS.n2150 VSS.t3405 11.0252
R9460 VSS.n2110 VSS.t4219 11.0252
R9461 VSS.n1893 VSS.t471 10.9418
R9462 VSS.n284 VSS.n283 10.5979
R9463 VSS.n2495 VSS.t58 10.5844
R9464 VSS.n2550 VSS.t336 10.5844
R9465 VSS.n1711 VSS.t791 10.5091
R9466 VSS.n1749 VSS.t2811 10.5091
R9467 VSS.n1916 VSS.t868 10.5091
R9468 VSS.n1992 VSS.t703 10.5091
R9469 VSS.n1340 VSS.t862 10.5091
R9470 VSS.n2029 VSS.t748 10.5091
R9471 VSS.n2039 VSS.t134 10.5091
R9472 VSS.n2045 VSS.t136 10.5091
R9473 VSS.n283 VSS.n282 10.4369
R9474 VSS.n281 VSS.n280 10.4308
R9475 VSS.n279 VSS.n278 10.4308
R9476 VSS.n277 VSS.n276 10.4308
R9477 VSS.n268 VSS.n266 10.357
R9478 VSS.n1708 VSS.t1720 10.2792
R9479 VSS.n1751 VSS.t2378 10.2792
R9480 VSS.n1912 VSS.t300 10.2792
R9481 VSS.n2021 VSS.t2691 10.2792
R9482 VSS.n1344 VSS.t4171 10.2792
R9483 VSS.n2026 VSS.t359 10.2792
R9484 VSS.n2036 VSS.t709 10.2792
R9485 VSS.n2047 VSS.t874 10.2792
R9486 VSS.n1700 VSS.t1730 10.2607
R9487 VSS.n1757 VSS.t2372 10.2607
R9488 VSS.n845 VSS.t304 10.2607
R9489 VSS.n2015 VSS.t2661 10.2607
R9490 VSS.n1353 VSS.t4169 10.2607
R9491 VSS.n743 VSS.t361 10.2607
R9492 VSS.n2031 VSS.t752 10.2607
R9493 VSS.n1345 VSS.t880 10.2607
R9494 VSS.n274 VSS.n273 10.2004
R9495 VSS.n270 VSS.n269 10.2004
R9496 VSS.n272 VSS.n271 10.198
R9497 VSS.n268 VSS.n267 10.1921
R9498 VSS.n524 VSS.t1794 9.93604
R9499 VSS.n1727 VSS.t2308 9.93604
R9500 VSS.n1729 VSS.t3792 9.93604
R9501 VSS.n1736 VSS.t2543 9.93604
R9502 VSS.n998 VSS.t2495 9.93604
R9503 VSS.n893 VSS.t841 9.93604
R9504 VSS.n1842 VSS.t1907 9.93604
R9505 VSS.n842 VSS.t902 9.93604
R9506 VSS.n2003 VSS.t4342 9.93604
R9507 VSS.n1991 VSS.t3805 9.93604
R9508 VSS.n1339 VSS.t3775 9.93604
R9509 VSS.n2043 VSS.t646 9.93604
R9510 VSS.n693 VSS.t4101 9.93604
R9511 VSS.n2062 VSS.t2415 9.93604
R9512 VSS.n2063 VSS.t3076 9.93604
R9513 VSS.n2003 VSS.t683 9.93029
R9514 VSS.n2117 VSS.t1110 9.93029
R9515 VSS.n1015 VSS.t4270 9.84591
R9516 VSS.n2096 VSS.t2875 9.84591
R9517 VSS.n2115 VSS.t3598 9.84591
R9518 VSS.n38 VSS.t379 9.84564
R9519 VSS.n19 VSS.t375 9.83796
R9520 VSS.n1978 VSS.t142 9.8287
R9521 VSS.n1966 VSS.t164 9.82208
R9522 VSS.n529 VSS.t3755 9.80518
R9523 VSS.n1017 VSS.t2319 9.80518
R9524 VSS.n976 VSS.t3699 9.80518
R9525 VSS.n918 VSS.t3433 9.80518
R9526 VSS.n930 VSS.t3321 9.80518
R9527 VSS.n894 VSS.t3683 9.80518
R9528 VSS.n895 VSS.t2614 9.80518
R9529 VSS.n860 VSS.t4035 9.80518
R9530 VSS.n874 VSS.t4148 9.80518
R9531 VSS.n869 VSS.t2521 9.80518
R9532 VSS.n791 VSS.t936 9.80518
R9533 VSS.n797 VSS.t3005 9.80518
R9534 VSS.n798 VSS.t1502 9.80518
R9535 VSS.n787 VSS.t1167 9.80518
R9536 VSS.n1998 VSS.t1905 9.80518
R9537 VSS.n753 VSS.t2951 9.80518
R9538 VSS.n1331 VSS.t1258 9.80518
R9539 VSS.n651 VSS.t4300 9.80518
R9540 VSS.n652 VSS.t2915 9.80518
R9541 VSS.n1453 VSS.t4291 9.80518
R9542 VSS.n417 VSS.t3163 9.80518
R9543 VSS.n421 VSS.t2196 9.80518
R9544 VSS.n1466 VSS.t2925 9.80518
R9545 VSS.n1462 VSS.t3956 9.80518
R9546 VSS.n1457 VSS.t2636 9.80518
R9547 VSS.n435 VSS.t1857 9.80518
R9548 VSS.n401 VSS.t435 9.80518
R9549 VSS.n1519 VSS.t2242 9.80518
R9550 VSS.n1513 VSS.t2343 9.80518
R9551 VSS.n617 VSS.t2407 9.80518
R9552 VSS.n609 VSS.t2417 9.80518
R9553 VSS.n605 VSS.t2481 9.80518
R9554 VSS.n626 VSS.t1510 9.80518
R9555 VSS.n1744 VSS.t3199 9.6277
R9556 VSS.n2040 VSS.t2802 9.6277
R9557 VSS.n742 VSS.t4181 9.6277
R9558 VSS.n2136 VSS.t1156 9.6277
R9559 VSS.n1833 VSS.t4226 9.38548
R9560 VSS.n1835 VSS.t4141 9.38548
R9561 VSS.n1210 VSS.t4134 9.38548
R9562 VSS.n852 VSS.t421 9.38548
R9563 VSS.n850 VSS.t4064 9.38548
R9564 VSS.n1913 VSS.t687 9.38548
R9565 VSS.n2151 VSS.t848 9.38548
R9566 VSS.n2149 VSS.t1129 9.38548
R9567 VSS.n38 VSS.t452 9.05755
R9568 VSS.n19 VSS.t462 9.05123
R9569 VSS.n18 VSS.n16 8.94121
R9570 VSS.n15 VSS.n13 8.94121
R9571 VSS.n44 VSS.n42 8.94121
R9572 VSS.n41 VSS.n39 8.94121
R9573 VSS.n923 VSS.t2539 8.63064
R9574 VSS.n907 VSS.t3157 8.63064
R9575 VSS.n866 VSS.t3376 8.63064
R9576 VSS.n718 VSS.t1203 8.63064
R9577 VSS.n2130 VSS.t4111 8.63064
R9578 VSS.n2214 VSS.t938 8.51132
R9579 VSS.n2247 VSS.t3781 8.51132
R9580 VSS.n2246 VSS.t1065 8.51132
R9581 VSS.n2245 VSS.t4230 8.51132
R9582 VSS.n2244 VSS.t3593 8.51132
R9583 VSS.n2243 VSS.t2399 8.51132
R9584 VSS.n2242 VSS.t3577 8.51132
R9585 VSS.n2241 VSS.t4119 8.51132
R9586 VSS.n2240 VSS.t4250 8.51132
R9587 VSS.n2238 VSS.t3292 8.51132
R9588 VSS.n2237 VSS.t1624 8.51132
R9589 VSS.n2236 VSS.t2341 8.51132
R9590 VSS.n2235 VSS.t2405 8.51132
R9591 VSS.n91 VSS.t4054 8.51132
R9592 VSS.n2315 VSS.t3803 8.51132
R9593 VSS.n2316 VSS.t2788 8.51132
R9594 VSS.n2317 VSS.t2465 8.51132
R9595 VSS.n2319 VSS.t3456 8.51132
R9596 VSS.n2320 VSS.t3379 8.51132
R9597 VSS.n2321 VSS.t3911 8.51132
R9598 VSS.n2322 VSS.t4175 8.51132
R9599 VSS.n2323 VSS.t3093 8.51132
R9600 VSS.n2324 VSS.t1522 8.51132
R9601 VSS.n2325 VSS.t2913 8.51132
R9602 VSS.n2326 VSS.t1524 8.51132
R9603 VSS.n2328 VSS.t3115 8.51132
R9604 VSS.n2327 VSS.t2054 8.51132
R9605 VSS.n89 VSS.t3801 8.51132
R9606 VSS.n2347 VSS.t1819 8.51132
R9607 VSS.n2346 VSS.t2325 8.51132
R9608 VSS.n2345 VSS.t2920 8.51132
R9609 VSS.n2344 VSS.t2136 8.51132
R9610 VSS.n2343 VSS.t3799 8.51132
R9611 VSS.n2341 VSS.t2621 8.51132
R9612 VSS.n2340 VSS.t2475 8.51132
R9613 VSS.n2339 VSS.t4327 8.51132
R9614 VSS.n2338 VSS.t3359 8.51132
R9615 VSS.n2337 VSS.t1583 8.51132
R9616 VSS.n2336 VSS.t1382 8.51132
R9617 VSS.n2335 VSS.t2850 8.51132
R9618 VSS.n2334 VSS.t4086 8.51132
R9619 VSS.n84 VSS.t4084 8.51132
R9620 VSS.n2408 VSS.t2089 8.51132
R9621 VSS.n2409 VSS.t3021 8.51132
R9622 VSS.n2410 VSS.t4082 8.51132
R9623 VSS.n2411 VSS.t3205 8.51132
R9624 VSS.n2413 VSS.t1734 8.51132
R9625 VSS.n2254 VSS.t2928 8.51132
R9626 VSS.n2256 VSS.t3905 8.51132
R9627 VSS.n2258 VSS.t1974 8.51132
R9628 VSS.n2260 VSS.t3037 8.51132
R9629 VSS.n2262 VSS.t3148 8.51132
R9630 VSS.n2264 VSS.t2885 8.51132
R9631 VSS.n2266 VSS.t4002 8.51132
R9632 VSS.n2280 VSS.t3934 8.51132
R9633 VSS.n2278 VSS.t2041 8.51132
R9634 VSS.n2276 VSS.t4329 8.51132
R9635 VSS.n2274 VSS.t3356 8.51132
R9636 VSS.n2272 VSS.t1247 8.51132
R9637 VSS.n2270 VSS.t3873 8.51132
R9638 VSS.n2268 VSS.t3526 8.51132
R9639 VSS.n2311 VSS.t2058 8.51132
R9640 VSS.n2309 VSS.t1184 8.51132
R9641 VSS.n2306 VSS.t2060 8.51132
R9642 VSS.n2304 VSS.t1186 8.51132
R9643 VSS.n2302 VSS.t2294 8.51132
R9644 VSS.n2300 VSS.t3207 8.51132
R9645 VSS.n2298 VSS.t3445 8.51132
R9646 VSS.n2296 VSS.t3250 8.51132
R9647 VSS.n2294 VSS.t1496 8.51132
R9648 VSS.n2292 VSS.t1874 8.51132
R9649 VSS.n2289 VSS.t3268 8.51132
R9650 VSS.n2287 VSS.t3907 8.51132
R9651 VSS.n2285 VSS.t3246 8.51132
R9652 VSS.n2283 VSS.t1301 8.51132
R9653 VSS.n87 VSS.t3861 8.51132
R9654 VSS.n2352 VSS.t4125 8.51132
R9655 VSS.n2354 VSS.t929 8.51132
R9656 VSS.n2356 VSS.t3855 8.51132
R9657 VSS.n2358 VSS.t2505 8.51132
R9658 VSS.n2361 VSS.t2549 8.51132
R9659 VSS.n2363 VSS.t1420 8.51132
R9660 VSS.n2365 VSS.t3427 8.51132
R9661 VSS.n2367 VSS.t3232 8.51132
R9662 VSS.n2369 VSS.t1233 8.51132
R9663 VSS.n2371 VSS.t2553 8.51132
R9664 VSS.n2373 VSS.t3256 8.51132
R9665 VSS.n2375 VSS.t3088 8.51132
R9666 VSS.n2380 VSS.t2585 8.51132
R9667 VSS.n2378 VSS.t1534 8.51132
R9668 VSS.n86 VSS.t3000 8.51132
R9669 VSS.n2402 VSS.t3211 8.51132
R9670 VSS.n2400 VSS.t3753 8.51132
R9671 VSS.n2398 VSS.t966 8.51132
R9672 VSS.n2396 VSS.t2536 8.51132
R9673 VSS.n2394 VSS.t974 8.51132
R9674 VSS.n2392 VSS.t2181 8.51132
R9675 VSS.n2389 VSS.t2638 8.51132
R9676 VSS.n2389 VSS.t3903 8.51132
R9677 VSS.n2388 VSS.t4132 8.51132
R9678 VSS.n2388 VSS.t3290 8.51132
R9679 VSS.n2387 VSS.t1943 8.51132
R9680 VSS.n2387 VSS.t3646 8.51132
R9681 VSS.n2386 VSS.t3313 8.51132
R9682 VSS.n2386 VSS.t2557 8.51132
R9683 VSS.n2385 VSS.t3013 8.51132
R9684 VSS.n2385 VSS.t3425 8.51132
R9685 VSS.n2384 VSS.t1455 8.51132
R9686 VSS.n2384 VSS.t1288 8.51132
R9687 VSS.n2383 VSS.t4155 8.51132
R9688 VSS.n2383 VSS.t2194 8.51132
R9689 VSS.n2382 VSS.t3518 8.51132
R9690 VSS.n2382 VSS.t1165 8.51132
R9691 VSS.n2390 VSS.t4096 8.51132
R9692 VSS.n2393 VSS.t1393 8.51132
R9693 VSS.n2395 VSS.t3123 8.51132
R9694 VSS.n2397 VSS.t3167 8.51132
R9695 VSS.n2399 VSS.t3230 8.51132
R9696 VSS.n2401 VSS.t3567 8.51132
R9697 VSS.n2403 VSS.t1030 8.51132
R9698 VSS.n2377 VSS.t1993 8.51132
R9699 VSS.n2379 VSS.t4129 8.51132
R9700 VSS.n2376 VSS.t3973 8.51132
R9701 VSS.n2374 VSS.t2492 8.51132
R9702 VSS.n2372 VSS.t1465 8.51132
R9703 VSS.n2370 VSS.t2140 8.51132
R9704 VSS.n2368 VSS.t1237 8.51132
R9705 VSS.n2366 VSS.t2247 8.51132
R9706 VSS.n2364 VSS.t3403 8.51132
R9707 VSS.n2362 VSS.t1461 8.51132
R9708 VSS.n2360 VSS.t4278 8.51132
R9709 VSS.n2357 VSS.t1758 8.51132
R9710 VSS.n2355 VSS.t2887 8.51132
R9711 VSS.n2353 VSS.t3409 8.51132
R9712 VSS.n2351 VSS.t3954 8.51132
R9713 VSS.n2282 VSS.t1506 8.51132
R9714 VSS.n2284 VSS.t3564 8.51132
R9715 VSS.n2286 VSS.t2168 8.51132
R9716 VSS.n2288 VSS.t1290 8.51132
R9717 VSS.n2291 VSS.t2033 8.51132
R9718 VSS.n2293 VSS.t1294 8.51132
R9719 VSS.n2295 VSS.t3150 8.51132
R9720 VSS.n2297 VSS.t2277 8.51132
R9721 VSS.n2299 VSS.t2111 8.51132
R9722 VSS.n2301 VSS.t1654 8.51132
R9723 VSS.n2303 VSS.t1708 8.51132
R9724 VSS.n2305 VSS.t2380 8.51132
R9725 VSS.n2307 VSS.t2228 8.51132
R9726 VSS.n2310 VSS.t1343 8.51132
R9727 VSS.n93 VSS.t2525 8.51132
R9728 VSS.n2269 VSS.t4341 8.51132
R9729 VSS.n2271 VSS.t2392 8.51132
R9730 VSS.n2273 VSS.t3896 8.51132
R9731 VSS.n2275 VSS.t1239 8.51132
R9732 VSS.n2277 VSS.t3511 8.51132
R9733 VSS.n2279 VSS.t3975 8.51132
R9734 VSS.n2267 VSS.t2455 8.51132
R9735 VSS.n2265 VSS.t3971 8.51132
R9736 VSS.n2263 VSS.t2652 8.51132
R9737 VSS.n2261 VSS.t3477 8.51132
R9738 VSS.n2259 VSS.t1699 8.51132
R9739 VSS.n2257 VSS.t978 8.51132
R9740 VSS.n2255 VSS.t3889 8.51132
R9741 VSS.n1143 VSS.t3487 8.51132
R9742 VSS.n1141 VSS.t3887 8.51132
R9743 VSS.n1139 VSS.t3727 8.51132
R9744 VSS.n1137 VSS.t4232 8.51132
R9745 VSS.n1135 VSS.t1262 8.51132
R9746 VSS.n1133 VSS.t1279 8.51132
R9747 VSS.n1131 VSS.t3190 8.51132
R9748 VSS.n1128 VSS.t2335 8.51132
R9749 VSS.n1126 VSS.t4252 8.51132
R9750 VSS.n1124 VSS.t1140 8.51132
R9751 VSS.n1122 VSS.t1474 8.51132
R9752 VSS.n1120 VSS.t955 8.51132
R9753 VSS.n1118 VSS.t2469 8.51132
R9754 VSS.n1116 VSS.t1001 8.51132
R9755 VSS.n1113 VSS.t1292 8.51132
R9756 VSS.n1111 VSS.t2234 8.51132
R9757 VSS.n1108 VSS.t1296 8.51132
R9758 VSS.n1106 VSS.t2287 8.51132
R9759 VSS.n1104 VSS.t1984 8.51132
R9760 VSS.n1102 VSS.t2828 8.51132
R9761 VSS.n1100 VSS.t3458 8.51132
R9762 VSS.n1098 VSS.t2771 8.51132
R9763 VSS.n1096 VSS.t2658 8.51132
R9764 VSS.n1094 VSS.t1587 8.51132
R9765 VSS.n1091 VSS.t4045 8.51132
R9766 VSS.n1089 VSS.t2605 8.51132
R9767 VSS.n1087 VSS.t2974 8.51132
R9768 VSS.n1085 VSS.t3925 8.51132
R9769 VSS.n1083 VSS.t957 8.51132
R9770 VSS.n1080 VSS.t3489 8.51132
R9771 VSS.n1078 VSS.t2608 8.51132
R9772 VSS.n1076 VSS.t2695 8.51132
R9773 VSS.n1074 VSS.t2836 8.51132
R9774 VSS.n1070 VSS.t1478 8.51132
R9775 VSS.n1068 VSS.t3892 8.51132
R9776 VSS.n1066 VSS.t2953 8.51132
R9777 VSS.n1064 VSS.t3626 8.51132
R9778 VSS.n1062 VSS.t3465 8.51132
R9779 VSS.n1060 VSS.t3763 8.51132
R9780 VSS.n1058 VSS.t1178 8.51132
R9781 VSS.n1056 VSS.t993 8.51132
R9782 VSS.n1054 VSS.t1090 8.51132
R9783 VSS.n1053 VSS.t2185 8.51132
R9784 VSS.n1053 VSS.t3357 8.51132
R9785 VSS.n1051 VSS.t1490 8.51132
R9786 VSS.n1051 VSS.t3806 8.51132
R9787 VSS.n1043 VSS.t948 8.51132
R9788 VSS.n1029 VSS.t3058 8.51132
R9789 VSS.n1031 VSS.t1695 8.51132
R9790 VSS.n1033 VSS.t3787 8.51132
R9791 VSS.n1035 VSS.t3656 8.51132
R9792 VSS.n1037 VSS.t2388 8.51132
R9793 VSS.n1039 VSS.t2224 8.51132
R9794 VSS.n1041 VSS.t1693 8.51132
R9795 VSS.n1044 VSS.t1669 8.51132
R9796 VSS.n1045 VSS.t3630 8.51132
R9797 VSS.n1047 VSS.t2261 8.51132
R9798 VSS.n1048 VSS.t997 8.51132
R9799 VSS.n1049 VSS.t4009 8.51132
R9800 VSS.n1050 VSS.t4335 8.51132
R9801 VSS.n1057 VSS.t2634 8.51132
R9802 VSS.n1059 VSS.t2347 8.51132
R9803 VSS.n1061 VSS.t2467 8.51132
R9804 VSS.n1063 VSS.t2962 8.51132
R9805 VSS.n1065 VSS.t2164 8.51132
R9806 VSS.n1067 VSS.t2555 8.51132
R9807 VSS.n1069 VSS.t2285 8.51132
R9808 VSS.n1071 VSS.t2354 8.51132
R9809 VSS.n1072 VSS.t4025 8.51132
R9810 VSS.n1075 VSS.t1152 8.51132
R9811 VSS.n1077 VSS.t3932 8.51132
R9812 VSS.n1079 VSS.t3286 8.51132
R9813 VSS.n1081 VSS.t3252 8.51132
R9814 VSS.n1084 VSS.t1716 8.51132
R9815 VSS.n1086 VSS.t2017 8.51132
R9816 VSS.n1088 VSS.t3936 8.51132
R9817 VSS.n1090 VSS.t2966 8.51132
R9818 VSS.n1093 VSS.t4019 8.51132
R9819 VSS.n1095 VSS.t2160 8.51132
R9820 VSS.n1097 VSS.t3452 8.51132
R9821 VSS.n1099 VSS.t1635 8.51132
R9822 VSS.n1101 VSS.t4217 8.51132
R9823 VSS.n1103 VSS.t3039 8.51132
R9824 VSS.n1105 VSS.t2901 8.51132
R9825 VSS.n1107 VSS.t2494 8.51132
R9826 VSS.n1109 VSS.t1551 8.51132
R9827 VSS.n1112 VSS.t1388 8.51132
R9828 VSS.n1115 VSS.t2323 8.51132
R9829 VSS.n1117 VSS.t1988 8.51132
R9830 VSS.n1119 VSS.t2958 8.51132
R9831 VSS.n1121 VSS.t1639 8.51132
R9832 VSS.n1123 VSS.t986 8.51132
R9833 VSS.n1125 VSS.t3033 8.51132
R9834 VSS.n1127 VSS.t2907 8.51132
R9835 VSS.n1130 VSS.t4322 8.51132
R9836 VSS.n1132 VSS.t3950 8.51132
R9837 VSS.n1134 VSS.t3101 8.51132
R9838 VSS.n1136 VSS.t1213 8.51132
R9839 VSS.n1138 VSS.t2899 8.51132
R9840 VSS.n1140 VSS.t3695 8.51132
R9841 VSS.n1142 VSS.t1530 8.51132
R9842 VSS.n1626 VSS.t2082 8.51132
R9843 VSS.n1628 VSS.t2289 8.51132
R9844 VSS.n1630 VSS.t1756 8.51132
R9845 VSS.n1632 VSS.t3390 8.51132
R9846 VSS.n1634 VSS.t1144 8.51132
R9847 VSS.n1636 VSS.t4152 8.51132
R9848 VSS.n1638 VSS.t2773 8.51132
R9849 VSS.n1641 VSS.t3960 8.51132
R9850 VSS.n1643 VSS.t3964 8.51132
R9851 VSS.n1645 VSS.t1919 8.51132
R9852 VSS.n1647 VSS.t4177 8.51132
R9853 VSS.n1649 VSS.t2064 8.51132
R9854 VSS.n1651 VSS.t1771 8.51132
R9855 VSS.n1653 VSS.t1406 8.51132
R9856 VSS.n1657 VSS.t3084 8.51132
R9857 VSS.n1659 VSS.t3713 8.51132
R9858 VSS.n1662 VSS.t3234 8.51132
R9859 VSS.n1664 VSS.t2070 8.51132
R9860 VSS.n1666 VSS.t2119 8.51132
R9861 VSS.n1668 VSS.t4242 8.51132
R9862 VSS.n1670 VSS.t1022 8.51132
R9863 VSS.n1672 VSS.t3562 8.51132
R9864 VSS.n1674 VSS.t4356 8.51132
R9865 VSS.n1676 VSS.t1375 8.51132
R9866 VSS.n1679 VSS.t3729 8.51132
R9867 VSS.n1681 VSS.t1034 8.51132
R9868 VSS.n1683 VSS.t4123 8.51132
R9869 VSS.n1685 VSS.t2463 8.51132
R9870 VSS.n1687 VSS.t1941 8.51132
R9871 VSS.n1690 VSS.t1915 8.51132
R9872 VSS.n1692 VSS.t1773 8.51132
R9873 VSS.n1694 VSS.t2479 8.51132
R9874 VSS.n1696 VSS.t4078 8.51132
R9875 VSS.n1723 VSS.t3788 8.51132
R9876 VSS.n1723 VSS.t1872 8.51132
R9877 VSS.n1722 VSS.t3450 8.51132
R9878 VSS.n1722 VSS.t3023 8.51132
R9879 VSS.n1721 VSS.t4127 8.51132
R9880 VSS.n1721 VSS.t4214 8.51132
R9881 VSS.n1720 VSS.t1746 8.51132
R9882 VSS.n1720 VSS.t2926 8.51132
R9883 VSS.n1724 VSS.t3041 8.51132
R9884 VSS.n1725 VSS.t2490 8.51132
R9885 VSS.n1733 VSS.t190 8.51132
R9886 VSS.n1713 VSS.t1235 8.51132
R9887 VSS.n1709 VSS.t991 8.51132
R9888 VSS.n1707 VSS.t4274 8.51132
R9889 VSS.n1705 VSS.t3176 8.51132
R9890 VSS.n1703 VSS.t2960 8.51132
R9891 VSS.n1701 VSS.t2598 8.51132
R9892 VSS.n1699 VSS.t2138 8.51132
R9893 VSS.n1698 VSS.t1243 8.51132
R9894 VSS.n1695 VSS.t2329 8.51132
R9895 VSS.n1693 VSS.t3182 8.51132
R9896 VSS.n1691 VSS.t3441 8.51132
R9897 VSS.n1689 VSS.t3520 8.51132
R9898 VSS.n1686 VSS.t1459 8.51132
R9899 VSS.n1684 VSS.t3485 8.51132
R9900 VSS.n1682 VSS.t3242 8.51132
R9901 VSS.n1680 VSS.t2595 8.51132
R9902 VSS.n1677 VSS.t2939 8.51132
R9903 VSS.n1675 VSS.t2786 8.51132
R9904 VSS.n1673 VSS.t1808 8.51132
R9905 VSS.n1671 VSS.t2964 8.51132
R9906 VSS.n1669 VSS.t3074 8.51132
R9907 VSS.n1667 VSS.t1764 8.51132
R9908 VSS.n1665 VSS.t2043 8.51132
R9909 VSS.n1663 VSS.t2712 8.51132
R9910 VSS.n1661 VSS.t4337 8.51132
R9911 VSS.n1658 VSS.t1227 8.51132
R9912 VSS.n1654 VSS.t2132 8.51132
R9913 VSS.n1652 VSS.t3339 8.51132
R9914 VSS.n1650 VSS.t1252 8.51132
R9915 VSS.n1648 VSS.t3019 8.51132
R9916 VSS.n1646 VSS.t1337 8.51132
R9917 VSS.n1644 VSS.t1853 8.51132
R9918 VSS.n1642 VSS.t3335 8.51132
R9919 VSS.n1639 VSS.t4276 8.51132
R9920 VSS.n1637 VSS.t3119 8.51132
R9921 VSS.n1635 VSS.t2212 8.51132
R9922 VSS.n1633 VSS.t3628 8.51132
R9923 VSS.n1631 VSS.t2183 8.51132
R9924 VSS.n1629 VSS.t2527 8.51132
R9925 VSS.n1627 VSS.t3551 8.51132
R9926 VSS.n1619 VSS.t3126 8.51132
R9927 VSS.n1617 VSS.t3555 8.51132
R9928 VSS.n1615 VSS.t2236 8.51132
R9929 VSS.n1613 VSS.t2449 8.51132
R9930 VSS.n1611 VSS.t1215 8.51132
R9931 VSS.n1609 VSS.t3048 8.51132
R9932 VSS.n1607 VSS.t3192 8.51132
R9933 VSS.n1604 VSS.t2403 8.51132
R9934 VSS.n1602 VSS.t4240 8.51132
R9935 VSS.n1600 VSS.t953 8.51132
R9936 VSS.n1598 VSS.t3522 8.51132
R9937 VSS.n1596 VSS.t3650 8.51132
R9938 VSS.n1594 VSS.t2703 8.51132
R9939 VSS.n1592 VSS.t1003 8.51132
R9940 VSS.n1589 VSS.t1298 8.51132
R9941 VSS.n1587 VSS.t2259 8.51132
R9942 VSS.n1584 VSS.t1422 8.51132
R9943 VSS.n1582 VSS.t1254 8.51132
R9944 VSS.n1580 VSS.t3715 8.51132
R9945 VSS.n1578 VSS.t3616 8.51132
R9946 VSS.n1576 VSS.t3463 8.51132
R9947 VSS.n1574 VSS.t3673 8.51132
R9948 VSS.n1572 VSS.t2697 8.51132
R9949 VSS.n1570 VSS.t2509 8.51132
R9950 VSS.n1567 VSS.t2121 8.51132
R9951 VSS.n1566 VSS.t4282 8.51132
R9952 VSS.n1566 VSS.t4213 8.51132
R9953 VSS.n1565 VSS.t2856 8.51132
R9954 VSS.n1565 VSS.t2942 8.51132
R9955 VSS.n1564 VSS.t2249 8.51132
R9956 VSS.n1564 VSS.t3537 8.51132
R9957 VSS.n971 VSS.t3144 8.51132
R9958 VSS.n971 VSS.t1492 8.51132
R9959 VSS.n1763 VSS.t2774 8.51132
R9960 VSS.n1763 VSS.t1476 8.51132
R9961 VSS.n1762 VSS.t2257 8.51132
R9962 VSS.n1762 VSS.t3890 8.51132
R9963 VSS.n1761 VSS.t4343 8.51132
R9964 VSS.n1761 VSS.t4154 8.51132
R9965 VSS.n1760 VSS.t2929 8.51132
R9966 VSS.n1760 VSS.t2832 8.51132
R9967 VSS.n993 VSS.t2056 8.51132
R9968 VSS.n995 VSS.t1273 8.51132
R9969 VSS.n1758 VSS.t1508 8.51132
R9970 VSS.n1569 VSS.t1245 8.51132
R9971 VSS.n1571 VSS.t3095 8.51132
R9972 VSS.n1573 VSS.t2541 8.51132
R9973 VSS.n1575 VSS.t3078 8.51132
R9974 VSS.n1577 VSS.t3794 8.51132
R9975 VSS.n1579 VSS.t3741 8.51132
R9976 VSS.n1581 VSS.t4298 8.51132
R9977 VSS.n1583 VSS.t2935 8.51132
R9978 VSS.n1585 VSS.t2830 8.51132
R9979 VSS.n1588 VSS.t2970 8.51132
R9980 VSS.n1591 VSS.t1882 8.51132
R9981 VSS.n1593 VSS.t3412 8.51132
R9982 VSS.n1595 VSS.t3418 8.51132
R9983 VSS.n1597 VSS.t3917 8.51132
R9984 VSS.n1599 VSS.t1775 8.51132
R9985 VSS.n1601 VSS.t2147 8.51132
R9986 VSS.n1603 VSS.t3325 8.51132
R9987 VSS.n1606 VSS.t2725 8.51132
R9988 VSS.n1608 VSS.t2871 8.51132
R9989 VSS.n1610 VSS.t3068 8.51132
R9990 VSS.n1612 VSS.t2972 8.51132
R9991 VSS.n1614 VSS.t4351 8.51132
R9992 VSS.n1616 VSS.t2721 8.51132
R9993 VSS.n1618 VSS.t2895 8.51132
R9994 VSS.n1176 VSS.t3503 8.51132
R9995 VSS.n1174 VSS.t4284 8.51132
R9996 VSS.n1172 VSS.t3509 8.51132
R9997 VSS.n1170 VSS.t2867 8.51132
R9998 VSS.n1168 VSS.t1615 8.51132
R9999 VSS.n1166 VSS.t961 8.51132
R10000 VSS.n1164 VSS.t4288 8.51132
R10001 VSS.n1161 VSS.t3844 8.51132
R10002 VSS.n1159 VSS.t1706 8.51132
R10003 VSS.n1157 VSS.t3044 8.51132
R10004 VSS.n1155 VSS.t2511 8.51132
R10005 VSS.n1153 VSS.t1482 8.51132
R10006 VSS.n1151 VSS.t1609 8.51132
R10007 VSS.n1149 VSS.t3645 8.51132
R10008 VSS.n1798 VSS.t3244 8.51132
R10009 VSS.n1796 VSS.t2166 8.51132
R10010 VSS.n1792 VSS.t2283 8.51132
R10011 VSS.n1790 VSS.t980 8.51132
R10012 VSS.n1788 VSS.t1965 8.51132
R10013 VSS.n1786 VSS.t3178 8.51132
R10014 VSS.n1784 VSS.t2158 8.51132
R10015 VSS.n1782 VSS.t3146 8.51132
R10016 VSS.n1780 VSS.t1028 8.51132
R10017 VSS.n1778 VSS.t3312 8.51132
R10018 VSS.n1776 VSS.t3539 8.51132
R10019 VSS.n1774 VSS.t1457 8.51132
R10020 VSS.n1772 VSS.t1864 8.51132
R10021 VSS.n1770 VSS.t1538 8.51132
R10022 VSS.n1768 VSS.t2854 8.51132
R10023 VSS.n968 VSS.t2386 8.51132
R10024 VSS.n967 VSS.t2006 8.51132
R10025 VSS.n957 VSS.t3443 8.51132
R10026 VSS.n969 VSS.t2707 8.51132
R10027 VSS.n1769 VSS.t3345 8.51132
R10028 VSS.n1771 VSS.t2798 8.51132
R10029 VSS.n1773 VSS.t2349 8.51132
R10030 VSS.n1775 VSS.t2411 8.51132
R10031 VSS.n1779 VSS.t4121 8.51132
R10032 VSS.n1781 VSS.t1589 8.51132
R10033 VSS.n1783 VSS.t3553 8.51132
R10034 VSS.n1785 VSS.t2019 8.51132
R10035 VSS.n1787 VSS.t3835 8.51132
R10036 VSS.n1789 VSS.t2547 8.51132
R10037 VSS.n1791 VSS.t4052 8.51132
R10038 VSS.n1793 VSS.t1884 8.51132
R10039 VSS.n1794 VSS.t968 8.51132
R10040 VSS.n1797 VSS.t2632 8.51132
R10041 VSS.n911 VSS.t3842 8.51132
R10042 VSS.n1150 VSS.t3534 8.51132
R10043 VSS.n1152 VSS.t1549 8.51132
R10044 VSS.n1154 VSS.t3624 8.51132
R10045 VSS.n1156 VSS.t2201 8.51132
R10046 VSS.n1158 VSS.t3665 8.51132
R10047 VSS.n1160 VSS.t2203 8.51132
R10048 VSS.n1163 VSS.t1652 8.51132
R10049 VSS.n1165 VSS.t3751 8.51132
R10050 VSS.n1167 VSS.t2623 8.51132
R10051 VSS.n1169 VSS.t1032 8.51132
R10052 VSS.n1171 VSS.t4006 8.51132
R10053 VSS.n1173 VSS.t1516 8.51132
R10054 VSS.n1175 VSS.t1591 8.51132
R10055 VSS.n1206 VSS.t3060 8.51132
R10056 VSS.n1204 VSS.t1760 8.51132
R10057 VSS.n1202 VSS.t2804 8.51132
R10058 VSS.n1200 VSS.t3507 8.51132
R10059 VSS.n1198 VSS.t3273 8.51132
R10060 VSS.n1196 VSS.t2729 8.51132
R10061 VSS.n1194 VSS.t1201 8.51132
R10062 VSS.n1191 VSS.t3254 8.51132
R10063 VSS.n1189 VSS.t3015 8.51132
R10064 VSS.n1187 VSS.t2699 8.51132
R10065 VSS.n1185 VSS.t2731 8.51132
R10066 VSS.n1183 VSS.t4029 8.51132
R10067 VSS.n1181 VSS.t4017 8.51132
R10068 VSS.n1179 VSS.t4173 8.51132
R10069 VSS.n1803 VSS.t2570 8.51132
R10070 VSS.n1805 VSS.t3765 8.51132
R10071 VSS.n1808 VSS.t2351 8.51132
R10072 VSS.n1810 VSS.t2834 8.51132
R10073 VSS.n1812 VSS.t3460 8.51132
R10074 VSS.n1814 VSS.t2937 8.51132
R10075 VSS.n1816 VSS.t2360 8.51132
R10076 VSS.n1818 VSS.t2778 8.51132
R10077 VSS.n1820 VSS.t4094 8.51132
R10078 VSS.n1822 VSS.t4011 8.51132
R10079 VSS.n1825 VSS.t3288 8.51132
R10080 VSS.n1827 VSS.t976 8.51132
R10081 VSS.n1830 VSS.t3240 8.51132
R10082 VSS.n1829 VSS.t2066 8.51132
R10083 VSS.n1828 VSS.t3454 8.51132
R10084 VSS.n1826 VSS.t2103 8.51132
R10085 VSS.n1823 VSS.t2903 8.51132
R10086 VSS.n1821 VSS.t2852 8.51132
R10087 VSS.n1819 VSS.t2149 8.51132
R10088 VSS.n1817 VSS.t3236 8.51132
R10089 VSS.n1815 VSS.t2390 8.51132
R10090 VSS.n1813 VSS.t2784 8.51132
R10091 VSS.n1811 VSS.t4302 8.51132
R10092 VSS.n1809 VSS.t3851 8.51132
R10093 VSS.n1807 VSS.t2956 8.51132
R10094 VSS.n1804 VSS.t3327 8.51132
R10095 VSS.n909 VSS.t3711 8.51132
R10096 VSS.n1180 VSS.t3885 8.51132
R10097 VSS.n1182 VSS.t4070 8.51132
R10098 VSS.n1184 VSS.t1663 8.51132
R10099 VSS.n1186 VSS.t2909 8.51132
R10100 VSS.n1188 VSS.t3394 8.51132
R10101 VSS.n1190 VSS.t4023 8.51132
R10102 VSS.n1193 VSS.t3025 8.51132
R10103 VSS.n1195 VSS.t3583 8.51132
R10104 VSS.n1197 VSS.t4244 8.51132
R10105 VSS.n1199 VSS.t3620 8.51132
R10106 VSS.n1201 VSS.t3154 8.51132
R10107 VSS.n1203 VSS.t1180 8.51132
R10108 VSS.n1205 VSS.t3679 8.51132
R10109 VSS.n1266 VSS.t3398 8.51132
R10110 VSS.n1264 VSS.t3938 8.51132
R10111 VSS.n1262 VSS.t1397 8.51132
R10112 VSS.n1260 VSS.t4345 8.51132
R10113 VSS.n1258 VSS.t1545 8.51132
R10114 VSS.n1256 VSS.t3228 8.51132
R10115 VSS.n1254 VSS.t2858 8.51132
R10116 VSS.n1251 VSS.t2445 8.51132
R10117 VSS.n1249 VSS.t3618 8.51132
R10118 VSS.n1247 VSS.t2737 8.51132
R10119 VSS.n1245 VSS.t3238 8.51132
R10120 VSS.n1243 VSS.t1917 8.51132
R10121 VSS.n1241 VSS.t3090 8.51132
R10122 VSS.n1239 VSS.t1468 8.51132
R10123 VSS.n1236 VSS.t2719 8.51132
R10124 VSS.n1234 VSS.t3827 8.51132
R10125 VSS.n1231 VSS.t2205 8.51132
R10126 VSS.n1229 VSS.t2616 8.51132
R10127 VSS.n1227 VSS.t3723 8.51132
R10128 VSS.n1225 VSS.t3350 8.51132
R10129 VSS.n1223 VSS.t3966 8.51132
R10130 VSS.n1221 VSS.t4272 8.51132
R10131 VSS.n1219 VSS.t3469 8.51132
R10132 VSS.n1217 VSS.t2877 8.51132
R10133 VSS.n1214 VSS.t2356 8.51132
R10134 VSS.n1213 VSS.t3671 8.51132
R10135 VSS.n886 VSS.t2230 8.51132
R10136 VSS.n1216 VSS.t1894 8.51132
R10137 VSS.n1218 VSS.t3305 8.51132
R10138 VSS.n1220 VSS.t4068 8.51132
R10139 VSS.n1222 VSS.t3103 8.51132
R10140 VSS.n1224 VSS.t2176 8.51132
R10141 VSS.n1226 VSS.t3923 8.51132
R10142 VSS.n1228 VSS.t3661 8.51132
R10143 VSS.n1230 VSS.t1886 8.51132
R10144 VSS.n1232 VSS.t1424 8.51132
R10145 VSS.n1235 VSS.t3364 8.51132
R10146 VSS.n1238 VSS.t1282 8.51132
R10147 VSS.n1240 VSS.t3303 8.51132
R10148 VSS.n1242 VSS.t1540 8.51132
R10149 VSS.n1244 VSS.t2333 8.51132
R10150 VSS.n1246 VSS.t2331 8.51132
R10151 VSS.n1248 VSS.t1714 8.51132
R10152 VSS.n1250 VSS.t3161 8.51132
R10153 VSS.n1253 VSS.t3224 8.51132
R10154 VSS.n1255 VSS.t3354 8.51132
R10155 VSS.n1257 VSS.t1649 8.51132
R10156 VSS.n1259 VSS.t1146 8.51132
R10157 VSS.n1261 VSS.t2933 8.51132
R10158 VSS.n1263 VSS.t2883 8.51132
R10159 VSS.n1265 VSS.t3818 8.51132
R10160 VSS.n1296 VSS.t2593 8.51132
R10161 VSS.n1294 VSS.t2382 8.51132
R10162 VSS.n1292 VSS.t4333 8.51132
R10163 VSS.n1290 VSS.t3424 8.51132
R10164 VSS.n1288 VSS.t3143 8.51132
R10165 VSS.n1286 VSS.t3536 8.51132
R10166 VSS.n1284 VSS.t1470 8.51132
R10167 VSS.n1281 VSS.t1020 8.51132
R10168 VSS.n1279 VSS.t1500 8.51132
R10169 VSS.n1277 VSS.t1931 8.51132
R10170 VSS.n1275 VSS.t3265 8.51132
R10171 VSS.n1273 VSS.t2447 8.51132
R10172 VSS.n1271 VSS.t4179 8.51132
R10173 VSS.n1269 VSS.t3602 8.51132
R10174 VSS.n1941 VSS.t1921 8.51132
R10175 VSS.n1939 VSS.t3894 8.51132
R10176 VSS.n1935 VSS.t2727 8.51132
R10177 VSS.n1933 VSS.t2897 8.51132
R10178 VSS.n1931 VSS.t2941 8.51132
R10179 VSS.n1929 VSS.t4150 8.51132
R10180 VSS.n1927 VSS.t1137 8.51132
R10181 VSS.n1925 VSS.t2705 8.51132
R10182 VSS.n1923 VSS.t1284 8.51132
R10183 VSS.n1921 VSS.t4144 8.51132
R10184 VSS.n1919 VSS.t1480 8.51132
R10185 VSS.n1917 VSS.t2485 8.51132
R10186 VSS.n1922 VSS.t3392 8.51132
R10187 VSS.n1924 VSS.t2645 8.51132
R10188 VSS.n1926 VSS.t1667 8.51132
R10189 VSS.n1928 VSS.t1617 8.51132
R10190 VSS.n1930 VSS.t1410 8.51132
R10191 VSS.n1932 VSS.t3881 8.51132
R10192 VSS.n1934 VSS.t2626 8.51132
R10193 VSS.n1936 VSS.t3731 8.51132
R10194 VSS.n1937 VSS.t1426 8.51132
R10195 VSS.n1940 VSS.t4146 8.51132
R10196 VSS.n780 VSS.t3226 8.51132
R10197 VSS.n1270 VSS.t2457 8.51132
R10198 VSS.n1272 VSS.t1327 8.51132
R10199 VSS.n1274 VSS.t3186 8.51132
R10200 VSS.n1276 VSS.t4258 8.51132
R10201 VSS.n1278 VSS.t3086 8.51132
R10202 VSS.n1280 VSS.t2419 8.51132
R10203 VSS.n1283 VSS.t3663 8.51132
R10204 VSS.n1285 VSS.t1339 8.51132
R10205 VSS.n1287 VSS.t3414 8.51132
R10206 VSS.n1289 VSS.t4280 8.51132
R10207 VSS.n1291 VSS.t2101 8.51132
R10208 VSS.n1293 VSS.t2198 8.51132
R10209 VSS.n1295 VSS.t3833 8.51132
R10210 VSS.n1326 VSS.t4354 8.51132
R10211 VSS.n1324 VSS.t2893 8.51132
R10212 VSS.n1322 VSS.t4339 8.51132
R10213 VSS.n1320 VSS.t1135 8.51132
R10214 VSS.n1318 VSS.t2086 8.51132
R10215 VSS.n1316 VSS.t2529 8.51132
R10216 VSS.n1314 VSS.t2487 8.51132
R10217 VSS.n1311 VSS.t3081 8.51132
R10218 VSS.n1309 VSS.t3174 8.51132
R10219 VSS.n1307 VSS.t3968 8.51132
R10220 VSS.n1305 VSS.t4228 8.51132
R10221 VSS.n1303 VSS.t3218 8.51132
R10222 VSS.n1301 VSS.t2507 8.51132
R10223 VSS.n1299 VSS.t1190 8.51132
R10224 VSS.n1946 VSS.t2619 8.51132
R10225 VSS.n1948 VSS.t2117 8.51132
R10226 VSS.n1952 VSS.t2848 8.51132
R10227 VSS.n1954 VSS.t2265 8.51132
R10228 VSS.n1956 VSS.t2358 8.51132
R10229 VSS.n1964 VSS.t4076 8.51132
R10230 VSS.n1962 VSS.t3869 8.51132
R10231 VSS.n1960 VSS.t1150 8.51132
R10232 VSS.n1958 VSS.t1211 8.51132
R10233 VSS.n1957 VSS.t3209 8.51132
R10234 VSS.n1955 VSS.t4234 8.51132
R10235 VSS.n1953 VSS.t4238 8.51132
R10236 VSS.n1951 VSS.t2780 8.51132
R10237 VSS.n1950 VSS.t4256 8.51132
R10238 VSS.n1947 VSS.t3808 8.51132
R10239 VSS.n778 VSS.t3479 8.51132
R10240 VSS.n1300 VSS.t3017 8.51132
R10241 VSS.n1302 VSS.t2409 8.51132
R10242 VSS.n1304 VSS.t3940 8.51132
R10243 VSS.n1306 VSS.t2072 8.51132
R10244 VSS.n1308 VSS.t3275 8.51132
R10245 VSS.n1310 VSS.t2968 8.51132
R10246 VSS.n1313 VSS.t2001 8.51132
R10247 VSS.n1315 VSS.t4021 8.51132
R10248 VSS.n1317 VSS.t1498 8.51132
R10249 VSS.n1319 VSS.t1395 8.51132
R10250 VSS.n1321 VSS.t2105 8.51132
R10251 VSS.n1323 VSS.t2985 8.51132
R10252 VSS.n1325 VSS.t2240 8.51132
R10253 VSS.n1397 VSS.t1892 8.51132
R10254 VSS.n1395 VSS.t1611 8.51132
R10255 VSS.n1393 VSS.t2483 8.51132
R10256 VSS.n1391 VSS.t2210 8.51132
R10257 VSS.n1389 VSS.t2820 8.51132
R10258 VSS.n1387 VSS.t2068 8.51132
R10259 VSS.n1385 VSS.t3783 8.51132
R10260 VSS.n1382 VSS.t2192 8.51132
R10261 VSS.n1381 VSS.t1567 8.51132
R10262 VSS.n1379 VSS.t1986 8.51132
R10263 VSS.n1377 VSS.t2782 8.51132
R10264 VSS.n1375 VSS.t3930 8.51132
R10265 VSS.n1373 VSS.t2327 8.51132
R10266 VSS.n1371 VSS.t1494 8.51132
R10267 VSS.n1368 VSS.t3248 8.51132
R10268 VSS.n1366 VSS.t3263 8.51132
R10269 VSS.n1362 VSS.t2564 8.51132
R10270 VSS.n1360 VSS.t1995 8.51132
R10271 VSS.n1358 VSS.t2568 8.51132
R10272 VSS.n1357 VSS.t2865 8.51132
R10273 VSS.n1355 VSS.t3366 8.51132
R10274 VSS.n1354 VSS.t4109 8.51132
R10275 VSS.n1350 VSS.t3825 8.51132
R10276 VSS.n1352 VSS.t1512 8.51132
R10277 VSS.n1361 VSS.t4027 8.51132
R10278 VSS.n1363 VSS.t2251 8.51132
R10279 VSS.n1364 VSS.t2987 8.51132
R10280 VSS.n1367 VSS.t1704 8.51132
R10281 VSS.n1370 VSS.t2701 8.51132
R10282 VSS.n1372 VSS.t2099 8.51132
R10283 VSS.n1374 VSS.t3333 8.51132
R10284 VSS.n1376 VSS.t3639 8.51132
R10285 VSS.n1378 VSS.t3652 8.51132
R10286 VSS.n1380 VSS.t4047 8.51132
R10287 VSS.n1384 VSS.t3216 8.51132
R10288 VSS.n1386 VSS.t3337 8.51132
R10289 VSS.n1388 VSS.t1659 8.51132
R10290 VSS.n1390 VSS.t4331 8.51132
R10291 VSS.n1392 VSS.t1444 8.51132
R10292 VSS.n1394 VSS.t1260 8.51132
R10293 VSS.n1396 VSS.t3871 8.51132
R10294 VSS.n1427 VSS.t4358 8.51132
R10295 VSS.n1425 VSS.t3258 8.51132
R10296 VSS.n1423 VSS.t3121 8.51132
R10297 VSS.n1421 VSS.t3913 8.51132
R10298 VSS.n1419 VSS.t3548 8.51132
R10299 VSS.n1417 VSS.t1665 8.51132
R10300 VSS.n1415 VSS.t2741 8.51132
R10301 VSS.n1412 VSS.t3180 8.51132
R10302 VSS.n1410 VSS.t3396 8.51132
R10303 VSS.n1408 VSS.t3952 8.51132
R10304 VSS.n1406 VSS.t1195 8.51132
R10305 VSS.n1404 VSS.t1963 8.51132
R10306 VSS.n1402 VSS.t3606 8.51132
R10307 VSS.n1400 VSS.t1225 8.51132
R10308 VSS.n2076 VSS.t3165 8.51132
R10309 VSS.n2074 VSS.t4066 8.51132
R10310 VSS.n2070 VSS.t2979 8.51132
R10311 VSS.n2068 VSS.t4131 8.51132
R10312 VSS.n2066 VSS.t2238 8.51132
R10313 VSS.n2065 VSS.t2869 8.51132
R10314 VSS.n2067 VSS.t4072 8.51132
R10315 VSS.n2069 VSS.t1241 8.51132
R10316 VSS.n2071 VSS.t2214 8.51132
R10317 VSS.n2072 VSS.t2654 8.51132
R10318 VSS.n2075 VSS.t1163 8.51132
R10319 VSS.n635 VSS.t1613 8.51132
R10320 VSS.n1401 VSS.t2142 8.51132
R10321 VSS.n1403 VSS.t2735 8.51132
R10322 VSS.n1405 VSS.t3996 8.51132
R10323 VSS.n1407 VSS.t3958 8.51132
R10324 VSS.n1409 VSS.t1565 8.51132
R10325 VSS.n1411 VSS.t2566 8.51132
R10326 VSS.n1414 VSS.t3921 8.51132
R10327 VSS.n1416 VSS.t3998 8.51132
R10328 VSS.n1418 VSS.t3648 8.51132
R10329 VSS.n1420 VSS.t2459 8.51132
R10330 VSS.n1422 VSS.t3613 8.51132
R10331 VSS.n1424 VSS.t3820 8.51132
R10332 VSS.n1426 VSS.t2226 8.51132
R10333 VSS.n1506 VSS.t2313 8.51132
R10334 VSS.n1504 VSS.t3481 8.51132
R10335 VSS.n1502 VSS.t1633 8.51132
R10336 VSS.n1500 VSS.t4056 8.51132
R10337 VSS.n1498 VSS.t972 8.51132
R10338 VSS.n1496 VSS.t3853 8.51132
R10339 VSS.n1494 VSS.t4347 8.51132
R10340 VSS.n1486 VSS.t3681 8.51132
R10341 VSS.n1484 VSS.t3416 8.51132
R10342 VSS.n1487 VSS.t2253 8.51132
R10343 VSS.n1490 VSS.t2009 8.51132
R10344 VSS.n1493 VSS.t2534 8.51132
R10345 VSS.n1495 VSS.t2113 8.51132
R10346 VSS.n1497 VSS.t2461 8.51132
R10347 VSS.n1499 VSS.t3611 8.51132
R10348 VSS.n1501 VSS.t4325 8.51132
R10349 VSS.n1503 VSS.t2413 8.51132
R10350 VSS.n1505 VSS.t1182 8.51132
R10351 VSS.n1528 VSS.t2640 8.51132
R10352 VSS.n1525 VSS.t3284 8.51132
R10353 VSS.n1529 VSS.t3188 8.51132
R10354 VSS.n1531 VSS.t2723 8.51132
R10355 VSS.n1539 VSS.t2097 8.51132
R10356 VSS.n1448 VSS.t2837 8.51132
R10357 VSS.n1448 VSS.t2717 8.51132
R10358 VSS.n1447 VSS.t3666 8.51132
R10359 VSS.n1447 VSS.t1142 8.51132
R10360 VSS.n1446 VSS.t4113 8.51132
R10361 VSS.n1446 VSS.t2232 8.51132
R10362 VSS.n1445 VSS.t1266 8.51132
R10363 VSS.n1445 VSS.t1552 8.51132
R10364 VSS.n1444 VSS.t1271 8.51132
R10365 VSS.n1444 VSS.t2278 8.51132
R10366 VSS.n1443 VSS.t1560 8.51132
R10367 VSS.n1443 VSS.t3116 8.51132
R10368 VSS.n1442 VSS.t4352 8.51132
R10369 VSS.n1442 VSS.t3294 8.51132
R10370 VSS.n1440 VSS.t1769 8.51132
R10371 VSS.n1439 VSS.t3821 8.51132
R10372 VSS.n1439 VSS.t3505 8.51132
R10373 VSS.n1438 VSS.t2401 8.51132
R10374 VSS.n1438 VSS.t3380 8.51132
R10375 VSS.n1437 VSS.t3857 8.51132
R10376 VSS.n1437 VSS.t3994 8.51132
R10377 VSS.n2082 VSS.t4211 8.51132
R10378 VSS.n2085 VSS.t2800 8.51132
R10379 VSS.n2083 VSS.t982 8.51132
R10380 VSS.n2081 VSS.t3384 8.51132
R10381 VSS.n1432 VSS.t1386 8.51132
R10382 VSS.n1433 VSS.t2739 8.51132
R10383 VSS.n1435 VSS.t1661 8.51132
R10384 VSS.n1888 VSS.t2513 8.49619
R10385 VSS.n834 VSS.t3172 8.49619
R10386 VSS.n699 VSS.t1080 8.47023
R10387 VSS.n697 VSS.t1078 8.47023
R10388 VSS.n1009 VSS.t3362 8.46241
R10389 VSS.n1014 VSS.t3675 8.46241
R10390 VSS.n933 VSS.t3725 8.46241
R10391 VSS.n1836 VSS.t2911 8.46241
R10392 VSS.n877 VSS.t2814 8.46241
R10393 VSS.n732 VSS.t2591 8.46241
R10394 VSS.n559 VSS.t3513 8.46241
R10395 VSS.n581 VSS.t465 8.46241
R10396 VSS.n2113 VSS.t2976 8.46241
R10397 VSS.n1986 VSS.t3139 8.44089
R10398 VSS.n1479 VSS.t3374 8.44089
R10399 VSS.n407 VSS.t1935 8.44089
R10400 VSS.n456 VSS.t3773 8.44089
R10401 VSS.n447 VSS.t4013 8.44089
R10402 VSS.n1436 VSS.t3879 8.44089
R10403 VSS.n690 VSS.t2123 8.43502
R10404 VSS.n692 VSS.t2126 8.43502
R10405 VSS.n1748 VSS.t2745 8.43208
R10406 VSS.n1010 VSS.t2889 8.43208
R10407 VSS.n945 VSS.t2130 8.43208
R10408 VSS.n940 VSS.t1645 8.43208
R10409 VSS.n958 VSS.t1710 8.43208
R10410 VSS.n1839 VSS.t4090 8.43208
R10411 VSS.n1875 VSS.t3769 8.43208
R10412 VSS.n884 VSS.t1038 8.43208
R10413 VSS.n1907 VSS.t1579 8.43208
R10414 VSS.n822 VSS.t1061 8.43208
R10415 VSS.n1990 VSS.t4039 8.43208
R10416 VSS.n2013 VSS.t3280 8.43208
R10417 VSS.n1984 VSS.t4246 8.43208
R10418 VSS.n738 VSS.t3029 8.43208
R10419 VSS.n2059 VSS.t1197 8.43208
R10420 VSS.n676 VSS.t1939 8.43208
R10421 VSS.n1474 VSS.t1903 8.43208
R10422 VSS.n560 VSS.t3431 8.43208
R10423 VSS.n562 VSS.t3632 8.43208
R10424 VSS.n2167 VSS.t3099 8.43208
R10425 VSS.n1526 VSS.t3499 8.43208
R10426 VSS.n441 VSS.t3735 8.43208
R10427 VSS.n444 VSS.t3689 8.43208
R10428 VSS.n455 VSS.t3515 8.43208
R10429 VSS.n2186 VSS.t3368 8.43208
R10430 VSS.n942 VSS.t1913 8.42575
R10431 VSS.n953 VSS.t1911 8.42575
R10432 VSS.n1876 VSS.t1909 8.42575
R10433 VSS.n1845 VSS.t1577 8.42575
R10434 VSS.n1887 VSS.t1131 8.42575
R10435 VSS.n831 VSS.t1878 8.42575
R10436 VSS.n733 VSS.t1311 8.42575
R10437 VSS.n686 VSS.t4183 8.42575
R10438 VSS.n687 VSS.t1949 8.42575
R10439 VSS.n596 VSS.t3220 8.42575
R10440 VSS.n2139 VSS.t1947 8.42575
R10441 VSS.n2142 VSS.t2747 8.42575
R10442 VSS.n2098 VSS.t3703 8.42575
R10443 VSS.n488 VSS.t3 8.4135
R10444 VSS.n1732 VSS.t4185 8.4135
R10445 VSS.n1735 VSS.t675 8.4135
R10446 VSS.n1013 VSS.t4196 8.4135
R10447 VSS.n1743 VSS.t2337 8.4135
R10448 VSS.n1747 VSS.t12 8.4135
R10449 VSS.n951 VSS.t2339 8.4135
R10450 VSS.n1212 VSS.t6 8.4135
R10451 VSS.n1915 VSS.t3902 8.4135
R10452 VSS.n1918 VSS.t4189 8.4135
R10453 VSS.n1970 VSS.t4193 8.4135
R10454 VSS.n2038 VSS.t3056 8.4135
R10455 VSS.n740 VSS.t1968 8.4135
R10456 VSS.n1346 VSS.t1074 8.4135
R10457 VSS.n2064 VSS.t1890 8.4135
R10458 VSS.n2061 VSS.t3697 8.4135
R10459 VSS.n675 VSS.t3309 8.4135
R10460 VSS.n597 VSS.t1123 8.4135
R10461 VSS.n446 VSS.t3307 8.4135
R10462 VSS.n2184 VSS.t3317 8.4135
R10463 VSS.n2138 VSS.t3677 8.4135
R10464 VSS.n2116 VSS.t834 8.4135
R10465 VSS.n2097 VSS.t2881 8.4135
R10466 VSS.n2086 VSS.t3319 8.4135
R10467 VSS.n833 VSS.t693 8.41154
R10468 VSS.n2048 VSS.t1117 8.41154
R10469 VSS.n944 VSS.t3296 8.4101
R10470 VSS.n956 VSS.t3737 8.4101
R10471 VSS.n1878 VSS.t1018 8.4101
R10472 VSS.n1843 VSS.t2503 8.4101
R10473 VSS.n1889 VSS.t2395 8.4101
R10474 VSS.n830 VSS.t2174 8.4101
R10475 VSS.n735 VSS.t995 8.4101
R10476 VSS.n689 VSS.t3323 8.4101
R10477 VSS.n685 VSS.t3105 8.4101
R10478 VSS.n2141 VSS.t2499 8.4101
R10479 VSS.n694 VSS.t1597 8.40958
R10480 VSS.n696 VSS.t1595 8.40958
R10481 VSS.n981 VSS.t2052 8.4005
R10482 VSS.n981 VSS.t515 8.4005
R10483 VSS.n986 VSS.t1005 8.4005
R10484 VSS.n986 VSS.t531 8.4005
R10485 VSS.n922 VSS.t499 8.4005
R10486 VSS.n922 VSS.t3072 8.4005
R10487 VSS.n931 VSS.t3875 8.4005
R10488 VSS.n931 VSS.t528 8.4005
R10489 VSS.n917 VSS.t488 8.4005
R10490 VSS.n917 VSS.t2153 8.4005
R10491 VSS.n902 VSS.t4107 8.4005
R10492 VSS.n902 VSS.t520 8.4005
R10493 VSS.n1856 VSS.t2317 8.4005
R10494 VSS.n1856 VSS.t510 8.4005
R10495 VSS.n875 VSS.t1133 8.4005
R10496 VSS.n875 VSS.t479 8.4005
R10497 VSS.n857 VSS.t4254 8.4005
R10498 VSS.n857 VSS.t780 8.4005
R10499 VSS.n805 VSS.t3757 8.4005
R10500 VSS.n805 VSS.t550 8.4005
R10501 VSS.n761 VSS.t490 8.4005
R10502 VSS.n761 VSS.t1536 8.4005
R10503 VSS.n1999 VSS.t1558 8.4005
R10504 VSS.n1999 VSS.t548 8.4005
R10505 VSS.n765 VSS.t814 8.4005
R10506 VSS.n765 VSS.t1256 8.4005
R10507 VSS.n727 VSS.t1063 8.4005
R10508 VSS.n727 VSS.t552 8.4005
R10509 VSS.n641 VSS.t1866 8.4005
R10510 VSS.n641 VSS.t778 8.4005
R10511 VSS.n659 VSS.t3046 8.4005
R10512 VSS.n659 VSS.t518 8.4005
R10513 VSS.n642 VSS.t830 8.4005
R10514 VSS.n642 VSS.t3035 8.4005
R10515 VSS.n1465 VSS.t3062 8.4005
R10516 VSS.n1465 VSS.t776 8.4005
R10517 VSS.n555 VSS.t774 8.4005
R10518 VSS.n555 VSS.t3596 8.4005
R10519 VSS.n547 VSS.t3009 8.4005
R10520 VSS.n547 VSS.t554 8.4005
R10521 VSS.n416 VSS.t3739 8.4005
R10522 VSS.n416 VSS.t546 8.4005
R10523 VSS.n1520 VSS.t1810 8.4005
R10524 VSS.n1520 VSS.t798 8.4005
R10525 VSS.n393 VSS.t802 8.4005
R10526 VSS.n393 VSS.t964 8.4005
R10527 VSS.n402 VSS.t782 8.4005
R10528 VSS.n402 VSS.t4004 8.4005
R10529 VSS.n433 VSS.t3654 8.4005
R10530 VSS.n433 VSS.t822 8.4005
R10531 VSS.n427 VSS.t2983 8.4005
R10532 VSS.n427 VSS.t824 8.4005
R10533 VSS.n616 VSS.t2049 8.4005
R10534 VSS.n616 VSS.t786 8.4005
R10535 VSS.n539 VSS.t2427 8.37615
R10536 VSS.n533 VSS.t2421 8.37615
R10537 VSS.n523 VSS.t2796 8.37615
R10538 VSS.n517 VSS.t3991 8.37615
R10539 VSS.n514 VSS.t1174 8.37615
R10540 VSS.n501 VSS.t451 8.37615
R10541 VSS.n497 VSS.t1742 8.37615
R10542 VSS.n491 VSS.t1785 8.37615
R10543 VSS.n487 VSS.t3131 8.37615
R10544 VSS.n2205 VSS.t1432 8.37615
R10545 VSS.n2207 VSS.t2574 8.37615
R10546 VSS.n2213 VSS.t236 8.37615
R10547 VSS.n2414 VSS.t942 8.37615
R10548 VSS.n2420 VSS.t699 8.37615
R10549 VSS.n1042 VSS.t4306 8.37615
R10550 VSS.n1030 VSS.t1053 8.37615
R10551 VSS.n1004 VSS.t3816 8.37615
R10552 VSS.n994 VSS.t1601 8.37615
R10553 VSS.n1871 VSS.t1750 8.37615
R10554 VSS.n1862 VSS.t314 8.37615
R10555 VSS.n1903 VSS.t1088 8.37615
R10556 VSS.n820 VSS.t1217 8.37615
R10557 VSS.n810 VSS.t53 8.37615
R10558 VSS.n839 VSS.t3759 8.37615
R10559 VSS.n674 VSS.t2995 8.37615
R10560 VSS.n664 VSS.t912 8.37615
R10561 VSS.n2164 VSS.t1446 8.37615
R10562 VSS.n564 VSS.t3747 8.37615
R10563 VSS.n574 VSS.t1675 8.37615
R10564 VSS.n2171 VSS.t1321 8.37615
R10565 VSS.n1540 VSS.t33 8.37615
R10566 VSS.n1530 VSS.t925 8.37615
R10567 VSS.n2193 VSS.t178 8.37615
R10568 VSS.n2185 VSS.t4262 8.37615
R10569 VSS.n590 VSS.t3495 8.37615
R10570 VSS.n580 VSS.t556 8.37615
R10571 VSS.n603 VSS.t3343 8.37615
R10572 VSS.n2102 VSS.t3709 8.36988
R10573 VSS.n1896 VSS.t468 8.3563
R10574 VSS.n836 VSS.t677 8.3563
R10575 VSS.n2044 VSS.t1112 8.3563
R10576 VSS.n18 VSS.n17 8.15207
R10577 VSS.n15 VSS.n14 8.15207
R10578 VSS.n44 VSS.n43 8.15207
R10579 VSS.n41 VSS.n40 8.15207
R10580 VSS.n2505 VSS.t339 7.60253
R10581 VSS.n29 VSS.t345 7.60253
R10582 VSS.n428 VSS.t3222 7.46717
R10583 VSS.n2127 VSS.t2749 7.46717
R10584 VSS.n2520 VSS.n2519 7.4193
R10585 VSS.n979 VSS.t534 7.3505
R10586 VSS.n983 VSS.t512 7.3505
R10587 VSS.n924 VSS.t522 7.3505
R10588 VSS.n929 VSS.t483 7.3505
R10589 VSS.n919 VSS.t524 7.3505
R10590 VSS.n903 VSS.t503 7.3505
R10591 VSS.n1854 VSS.t485 7.3505
R10592 VSS.n873 VSS.t506 7.3505
R10593 VSS.n854 VSS.t790 7.3505
R10594 VSS.n802 VSS.t495 7.3505
R10595 VSS.n759 VSS.t538 7.3505
R10596 VSS.n1997 VSS.t492 7.3505
R10597 VSS.n762 VSS.t811 7.3505
R10598 VSS.n726 VSS.t497 7.3505
R10599 VSS.n638 VSS.t784 7.3505
R10600 VSS.n656 VSS.t536 7.3505
R10601 VSS.n645 VSS.t768 7.3505
R10602 VSS.n1463 VSS.t807 7.3505
R10603 VSS.n553 VSS.t764 7.3505
R10604 VSS.n550 VSS.t543 7.3505
R10605 VSS.n414 VSS.t481 7.3505
R10606 VSS.n1518 VSS.t809 7.3505
R10607 VSS.n438 VSS.t794 7.3505
R10608 VSS.n434 VSS.t828 7.3505
R10609 VSS.n424 VSS.t818 7.3505
R10610 VSS.n396 VSS.t766 7.3505
R10611 VSS.n618 VSS.t805 7.3505
R10612 VSS.n2533 VSS.n2532 7.344
R10613 VSS.n2518 VSS.n2517 7.25447
R10614 VSS.n2475 VSS.t192 7.21552
R10615 VSS.n119 VSS.t1924 7.21552
R10616 VSS.n148 VSS.t413 7.21552
R10617 VSS.n177 VSS.t65 7.21552
R10618 VSS.n206 VSS.t121 7.21552
R10619 VSS.n235 VSS.t565 7.21552
R10620 VSS.n290 VSS.t2759 7.21552
R10621 VSS.n326 VSS.t113 7.21552
R10622 VSS.n1712 VSS.t3201 7.06906
R10623 VSS.n623 VSS.t1071 7.06906
R10624 VSS.n610 VSS.t1563 7.06906
R10625 VSS.n29 VSS.t888 6.81584
R10626 VSS.n2505 VSS.t895 6.81584
R10627 VSS.n10 VSS.t1976 6.80897
R10628 VSS.n9 VSS.t417 6.80897
R10629 VSS.n8 VSS.t73 6.80897
R10630 VSS.n7 VSS.t125 6.80897
R10631 VSS.n6 VSS.t559 6.80897
R10632 VSS.t2766 VSS.n4 6.80897
R10633 VSS.n5 VSS.t105 6.80897
R10634 VSS.n2551 VSS.t196 6.80897
R10635 VSS.n2550 VSS.n10 6.73275
R10636 VSS.n2550 VSS.n9 6.73275
R10637 VSS.n2550 VSS.n8 6.73275
R10638 VSS.n2550 VSS.n7 6.73275
R10639 VSS.n2550 VSS.n6 6.73275
R10640 VSS.n2550 VSS.n4 6.73275
R10641 VSS.n2550 VSS.n5 6.73275
R10642 VSS.n2551 VSS.n2550 6.73275
R10643 VSS.n28 VSS.n26 6.70371
R10644 VSS.n25 VSS.n23 6.70371
R10645 VSS.n2501 VSS.n2499 6.70371
R10646 VSS.n2504 VSS.n2502 6.70371
R10647 VSS.n479 VSS.t4103 6.63343
R10648 VSS.n1718 VSS.t1378 6.63343
R10649 VSS.n914 VSS.t2393 6.63343
R10650 VSS.n864 VSS.t4060 6.63343
R10651 VSS.n1209 VSS.t4224 6.63343
R10652 VSS.n801 VSS.t900 6.63343
R10653 VSS.n460 VSS.t2269 6.63343
R10654 VSS.n630 VSS.t3544 6.63343
R10655 VSS.n629 VSS.t129 6.63343
R10656 VSS.n624 VSS.t1069 6.63343
R10657 VSS.n1746 VSS.n979 6.55876
R10658 VSS.n1008 VSS.n983 6.55876
R10659 VSS.n947 VSS.n924 6.55876
R10660 VSS.n938 VSS.n929 6.55876
R10661 VSS.n959 VSS.n919 6.55876
R10662 VSS.n1841 VSS.n903 6.55876
R10663 VSS.n1872 VSS.n1854 6.55876
R10664 VSS.n882 VSS.n873 6.55876
R10665 VSS.n1905 VSS.n854 6.55876
R10666 VSS.n819 VSS.n802 6.55876
R10667 VSS.n1988 VSS.n759 6.55876
R10668 VSS.n2010 VSS.n1997 6.55876
R10669 VSS.n1982 VSS.n762 6.55876
R10670 VSS.n736 VSS.n726 6.55876
R10671 VSS.n2057 VSS.n638 6.55876
R10672 VSS.n673 VSS.n656 6.55876
R10673 VSS.n698 VSS.n645 6.55876
R10674 VSS.n1473 VSS.n1463 6.55876
R10675 VSS.n558 VSS.n553 6.55876
R10676 VSS.n565 VSS.n550 6.55876
R10677 VSS.n2165 VSS.n414 6.55876
R10678 VSS.n1523 VSS.n1518 6.55876
R10679 VSS.n439 VSS.n438 6.55876
R10680 VSS.n445 VSS.n434 6.55876
R10681 VSS.n425 VSS.n424 6.55876
R10682 VSS.n2188 VSS.n396 6.55876
R10683 VSS.n2104 VSS.n618 6.55876
R10684 VSS.n2041 VSS.n709 6.52354
R10685 VSS.n1714 VSS.n1712 6.4805
R10686 VSS.n2094 VSS.n623 6.4805
R10687 VSS.n2114 VSS.n610 6.4805
R10688 VSS.n589 VSS.n461 6.47521
R10689 VSS.n2147 VSS.n606 6.47521
R10690 VSS.n584 VSS.n465 6.46859
R10691 VSS.n594 VSS.n428 6.46859
R10692 VSS.n2151 VSS.n604 6.46859
R10693 VSS.n2144 VSS.n2127 6.46859
R10694 VSS.n1011 VSS.n982 6.46615
R10695 VSS.n1000 VSS.n989 6.46615
R10696 VSS.n955 VSS.n920 6.46615
R10697 VSS.n934 VSS.n932 6.46615
R10698 VSS.n966 VSS.n913 6.46615
R10699 VSS.n1849 VSS.n899 6.46615
R10700 VSS.n1864 VSS.n1860 6.46615
R10701 VSS.n878 VSS.n876 6.46615
R10702 VSS.n1898 VSS.n859 6.46615
R10703 VSS.n811 VSS.n809 6.46615
R10704 VSS.n1981 VSS.n763 6.46615
R10705 VSS.n2005 VSS.n2001 6.46615
R10706 VSS.n1973 VSS.n769 6.46615
R10707 VSS.n730 VSS.n729 6.46615
R10708 VSS.n701 VSS.n643 6.46615
R10709 VSS.n665 VSS.n663 6.46615
R10710 VSS.n2055 VSS.n640 6.46615
R10711 VSS.n1468 VSS.n1467 6.46615
R10712 VSS.n2157 VSS.n420 6.46615
R10713 VSS.n573 VSS.n543 6.46615
R10714 VSS.n2159 VSS.n418 6.46615
R10715 VSS.n2197 VSS.n388 6.46615
R10716 VSS.n2181 VSS.n400 6.46615
R10717 VSS.n452 VSS.n430 6.46615
R10718 VSS.n593 VSS.n429 6.46615
R10719 VSS.n2196 VSS.n389 6.46615
R10720 VSS.n2111 VSS.n612 6.46615
R10721 VSS.n1710 VSS.n1019 6.46462
R10722 VSS.n1750 VSS.n978 6.46462
R10723 VSS.n1914 VSS.n782 6.46462
R10724 VSS.n1959 VSS.n777 6.46462
R10725 VSS.n1961 VSS.n776 6.46462
R10726 VSS.n1963 VSS.n775 6.46462
R10727 VSS.n751 VSS.n750 6.46462
R10728 VSS.n1342 VSS.n1337 6.46462
R10729 VSS.n2027 VSS.n717 6.46462
R10730 VSS.n2037 VSS.n710 6.46462
R10731 VSS.n2046 VSS.n707 6.46462
R10732 VSS.n1702 VSS.n1022 6.45138
R10733 VSS.n1704 VSS.n1021 6.45138
R10734 VSS.n1706 VSS.n1020 6.45138
R10735 VSS.n1752 VSS.n977 6.45138
R10736 VSS.n1754 VSS.n975 6.45138
R10737 VSS.n1755 VSS.n974 6.45138
R10738 VSS.n849 VSS.n783 6.45138
R10739 VSS.n848 VSS.n784 6.45138
R10740 VSS.n846 VSS.n786 6.45138
R10741 VSS.n1967 VSS.n773 6.45138
R10742 VSS.n1968 VSS.n772 6.45138
R10743 VSS.n1969 VSS.n771 6.45138
R10744 VSS.n1971 VSS.n770 6.45138
R10745 VSS.n1974 VSS.n768 6.45138
R10746 VSS.n1976 VSS.n767 6.45138
R10747 VSS.n1977 VSS.n766 6.45138
R10748 VSS.n2020 VSS.n752 6.45138
R10749 VSS.n2018 VSS.n754 6.45138
R10750 VSS.n2017 VSS.n755 6.45138
R10751 VSS.n1351 VSS.n1332 6.45138
R10752 VSS.n1348 VSS.n1334 6.45138
R10753 VSS.n1347 VSS.n1335 6.45138
R10754 VSS.n744 VSS.n722 6.45138
R10755 VSS.n746 VSS.n720 6.45138
R10756 VSS.n747 VSS.n719 6.45138
R10757 VSS.n2033 VSS.n713 6.45138
R10758 VSS.n2034 VSS.n712 6.45138
R10759 VSS.n2035 VSS.n711 6.45138
R10760 VSS.n706 VSS.n705 6.45138
R10761 VSS.n1341 VSS.n1338 6.45138
R10762 VSS.n1343 VSS.n1336 6.45138
R10763 VSS.n516 VSS.n479 6.45115
R10764 VSS.n1728 VSS.n1718 6.45115
R10765 VSS.n965 VSS.n914 6.45115
R10766 VSS.n1891 VSS.n864 6.45115
R10767 VSS.n1211 VSS.n1209 6.45115
R10768 VSS.n821 VSS.n801 6.45115
R10769 VSS.n591 VSS.n460 6.45115
R10770 VSS.n2087 VSS.n630 6.45115
R10771 VSS.n2088 VSS.n629 6.45115
R10772 VSS.n2093 VSS.n624 6.45115
R10773 VSS.n1989 VSS.n758 6.44333
R10774 VSS.n1987 VSS.n760 6.44333
R10775 VSS.n1478 VSS.n1459 6.44333
R10776 VSS.n1476 VSS.n1461 6.44333
R10777 VSS.n2173 VSS.n408 6.44333
R10778 VSS.n2170 VSS.n410 6.44333
R10779 VSS.n599 VSS.n426 6.44333
R10780 VSS.n454 VSS.n453 6.44333
R10781 VSS.n450 VSS.n431 6.44333
R10782 VSS.n449 VSS.n432 6.44333
R10783 VSS.n1434 VSS.n1431 6.44333
R10784 VSS.n633 VSS.n632 6.44333
R10785 VSS.n1742 VSS.n981 6.43285
R10786 VSS.n1005 VSS.n986 6.43285
R10787 VSS.n950 VSS.n922 6.43285
R10788 VSS.n936 VSS.n931 6.43285
R10789 VSS.n961 VSS.n917 6.43285
R10790 VSS.n1844 VSS.n902 6.43285
R10791 VSS.n1869 VSS.n1856 6.43285
R10792 VSS.n880 VSS.n875 6.43285
R10793 VSS.n1901 VSS.n857 6.43285
R10794 VSS.n816 VSS.n805 6.43285
R10795 VSS.n1985 VSS.n761 6.43285
R10796 VSS.n2008 VSS.n1999 6.43285
R10797 VSS.n1979 VSS.n765 6.43285
R10798 VSS.n734 VSS.n727 6.43285
R10799 VSS.n2054 VSS.n641 6.43285
R10800 VSS.n670 VSS.n659 6.43285
R10801 VSS.n702 VSS.n642 6.43285
R10802 VSS.n1471 VSS.n1465 6.43285
R10803 VSS.n556 VSS.n555 6.43285
R10804 VSS.n568 VSS.n547 6.43285
R10805 VSS.n2162 VSS.n416 6.43285
R10806 VSS.n1521 VSS.n1520 6.43285
R10807 VSS.n2191 VSS.n393 6.43285
R10808 VSS.n2178 VSS.n402 6.43285
R10809 VSS.n448 VSS.n433 6.43285
R10810 VSS.n598 VSS.n427 6.43285
R10811 VSS.n2106 VSS.n616 6.43285
R10812 VSS.n540 VSS.n468 6.41829
R10813 VSS.n502 VSS.n498 6.41829
R10814 VSS.n490 VSS.n485 6.41829
R10815 VSS.n2407 VSS.n83 6.41829
R10816 VSS.n1726 VSS.n1719 6.41829
R10817 VSS.n1731 VSS.n1018 6.41829
R10818 VSS.n1006 VSS.n985 6.41829
R10819 VSS.n1831 VSS.n908 6.41829
R10820 VSS.n1873 VSS.n1853 6.41829
R10821 VSS.n1877 VSS.n898 6.41829
R10822 VSS.n1906 VSS.n853 6.41829
R10823 VSS.n1895 VSS.n861 6.41829
R10824 VSS.n1892 VSS.n863 6.41829
R10825 VSS.n835 VSS.n793 6.41829
R10826 VSS.n824 VSS.n799 6.41829
R10827 VSS.n847 VSS.n785 6.41829
R10828 VSS.n2014 VSS.n757 6.41829
R10829 VSS.n2007 VSS.n2000 6.41829
R10830 VSS.n730 VSS.n728 6.41829
R10831 VSS.n683 VSS.n649 6.41829
R10832 VSS.n682 VSS.n650 6.41829
R10833 VSS.n2056 VSS.n639 6.41829
R10834 VSS.n2058 VSS.n637 6.41829
R10835 VSS.n1482 VSS.n1456 6.41829
R10836 VSS.n563 VSS.n551 6.41829
R10837 VSS.n1488 VSS.n1454 6.41829
R10838 VSS.n2183 VSS.n398 6.41829
R10839 VSS.n2090 VSS.n627 6.41829
R10840 VSS.n2092 VSS.n625 6.41829
R10841 VSS.n2099 VSS.n621 6.41829
R10842 VSS.n2101 VSS.n619 6.41829
R10843 VSS.n2112 VSS.n611 6.41829
R10844 VSS.n2135 VSS.n2131 6.41829
R10845 VSS.n2134 VSS.n2132 6.41829
R10846 VSS.n2004 VSS.n2002 6.40771
R10847 VSS.n2119 VSS.n608 6.40771
R10848 VSS.n1894 VSS.n862 6.39182
R10849 VSS.n530 VSS.n529 6.38659
R10850 VSS.n1734 VSS.n1017 6.38659
R10851 VSS.n1753 VSS.n976 6.38659
R10852 VSS.n960 VSS.n918 6.38659
R10853 VSS.n937 VSS.n930 6.38659
R10854 VSS.n948 VSS.n923 6.38659
R10855 VSS.n1882 VSS.n894 6.38659
R10856 VSS.n1881 VSS.n895 6.38659
R10857 VSS.n1834 VSS.n907 6.38659
R10858 VSS.n1897 VSS.n860 6.38659
R10859 VSS.n891 VSS.n866 6.38659
R10860 VSS.n881 VSS.n874 6.38659
R10861 VSS.n888 VSS.n869 6.38659
R10862 VSS.n838 VSS.n791 6.38659
R10863 VSS.n826 VSS.n797 6.38659
R10864 VSS.n825 VSS.n798 6.38659
R10865 VSS.n844 VSS.n787 6.38659
R10866 VSS.n2009 VSS.n1998 6.38659
R10867 VSS.n2019 VSS.n753 6.38659
R10868 VSS.n748 VSS.n718 6.38659
R10869 VSS.n1356 VSS.n1331 6.38659
R10870 VSS.n681 VSS.n651 6.38659
R10871 VSS.n680 VSS.n652 6.38659
R10872 VSS.n1489 VSS.n1453 6.38659
R10873 VSS.n2161 VSS.n417 6.38659
R10874 VSS.n422 VSS.n421 6.38659
R10875 VSS.n1469 VSS.n1466 6.38659
R10876 VSS.n1475 VSS.n1462 6.38659
R10877 VSS.n1481 VSS.n1457 6.38659
R10878 VSS.n443 VSS.n435 6.38659
R10879 VSS.n2179 VSS.n401 6.38659
R10880 VSS.n1522 VSS.n1519 6.38659
R10881 VSS.n1534 VSS.n1513 6.38659
R10882 VSS.n2105 VSS.n617 6.38659
R10883 VSS.n2118 VSS.n609 6.38659
R10884 VSS.n2148 VSS.n605 6.38659
R10885 VSS.n2137 VSS.n2130 6.38659
R10886 VSS.n2091 VSS.n626 6.38659
R10887 VSS.n1848 VSS.n900 6.38521
R10888 VSS.n1846 VSS.n901 6.38521
R10889 VSS.n538 VSS.n469 6.37859
R10890 VSS.n537 VSS.n470 6.37859
R10891 VSS.n536 VSS.n471 6.37859
R10892 VSS.n535 VSS.n472 6.37859
R10893 VSS.n534 VSS.n473 6.37859
R10894 VSS.n522 VSS.n474 6.37859
R10895 VSS.n521 VSS.n475 6.37859
R10896 VSS.n520 VSS.n476 6.37859
R10897 VSS.n519 VSS.n477 6.37859
R10898 VSS.n518 VSS.n478 6.37859
R10899 VSS.n513 VSS.n506 6.37859
R10900 VSS.n512 VSS.n507 6.37859
R10901 VSS.n511 VSS.n508 6.37859
R10902 VSS.n510 VSS.n509 6.37859
R10903 VSS.n500 VSS.n499 6.37859
R10904 VSS.n496 VSS.n480 6.37859
R10905 VSS.n495 VSS.n481 6.37859
R10906 VSS.n494 VSS.n482 6.37859
R10907 VSS.n493 VSS.n483 6.37859
R10908 VSS.n492 VSS.n484 6.37859
R10909 VSS.n385 VSS.n384 6.37859
R10910 VSS.n2201 VSS.n383 6.37859
R10911 VSS.n2202 VSS.n382 6.37859
R10912 VSS.n2203 VSS.n381 6.37859
R10913 VSS.n2204 VSS.n380 6.37859
R10914 VSS.n2208 VSS.n378 6.37859
R10915 VSS.n2209 VSS.n377 6.37859
R10916 VSS.n2210 VSS.n376 6.37859
R10917 VSS.n2211 VSS.n375 6.37859
R10918 VSS.n2212 VSS.n374 6.37859
R10919 VSS.n2415 VSS.n81 6.37859
R10920 VSS.n2416 VSS.n80 6.37859
R10921 VSS.n2417 VSS.n79 6.37859
R10922 VSS.n2418 VSS.n78 6.37859
R10923 VSS.n2419 VSS.n77 6.37859
R10924 VSS.n1040 VSS.n1024 6.37859
R10925 VSS.n1038 VSS.n1025 6.37859
R10926 VSS.n1036 VSS.n1026 6.37859
R10927 VSS.n1034 VSS.n1027 6.37859
R10928 VSS.n1032 VSS.n1028 6.37859
R10929 VSS.n1003 VSS.n987 6.37859
R10930 VSS.n1001 VSS.n988 6.37859
R10931 VSS.n999 VSS.n990 6.37859
R10932 VSS.n997 VSS.n991 6.37859
R10933 VSS.n996 VSS.n992 6.37859
R10934 VSS.n1870 VSS.n1855 6.37859
R10935 VSS.n1868 VSS.n1857 6.37859
R10936 VSS.n1867 VSS.n1858 6.37859
R10937 VSS.n1866 VSS.n1859 6.37859
R10938 VSS.n1863 VSS.n1861 6.37859
R10939 VSS.n1904 VSS.n855 6.37859
R10940 VSS.n818 VSS.n803 6.37859
R10941 VSS.n817 VSS.n804 6.37859
R10942 VSS.n815 VSS.n806 6.37859
R10943 VSS.n814 VSS.n807 6.37859
R10944 VSS.n812 VSS.n808 6.37859
R10945 VSS.n837 VSS.n792 6.37859
R10946 VSS.n672 VSS.n657 6.37859
R10947 VSS.n671 VSS.n658 6.37859
R10948 VSS.n669 VSS.n660 6.37859
R10949 VSS.n668 VSS.n661 6.37859
R10950 VSS.n666 VSS.n662 6.37859
R10951 VSS.n2166 VSS.n413 6.37859
R10952 VSS.n566 VSS.n549 6.37859
R10953 VSS.n567 VSS.n548 6.37859
R10954 VSS.n569 VSS.n546 6.37859
R10955 VSS.n570 VSS.n545 6.37859
R10956 VSS.n572 VSS.n544 6.37859
R10957 VSS.n2169 VSS.n411 6.37859
R10958 VSS.n1538 VSS.n1509 6.37859
R10959 VSS.n1536 VSS.n1511 6.37859
R10960 VSS.n1535 VSS.n1512 6.37859
R10961 VSS.n1533 VSS.n1514 6.37859
R10962 VSS.n1532 VSS.n1515 6.37859
R10963 VSS.n2192 VSS.n391 6.37859
R10964 VSS.n2191 VSS.n392 6.37859
R10965 VSS.n2190 VSS.n394 6.37859
R10966 VSS.n2189 VSS.n395 6.37859
R10967 VSS.n2187 VSS.n397 6.37859
R10968 VSS.n588 VSS.n462 6.37859
R10969 VSS.n587 VSS.n463 6.37859
R10970 VSS.n585 VSS.n464 6.37859
R10971 VSS.n583 VSS.n466 6.37859
R10972 VSS.n582 VSS.n467 6.37859
R10973 VSS.n2122 VSS.n2121 6.37859
R10974 VSS.n2100 VSS.n620 6.37859
R10975 VSS.n531 VSS.n528 6.35874
R10976 VSS.n1737 VSS.n1016 6.35874
R10977 VSS.n1756 VSS.n973 6.35874
R10978 VSS.n962 VSS.n916 6.35874
R10979 VSS.n939 VSS.n928 6.35874
R10980 VSS.n943 VSS.n926 6.35874
R10981 VSS.n946 VSS.n925 6.35874
R10982 VSS.n1880 VSS.n896 6.35874
R10983 VSS.n1879 VSS.n897 6.35874
R10984 VSS.n1840 VSS.n904 6.35874
R10985 VSS.n1837 VSS.n906 6.35874
R10986 VSS.n1900 VSS.n858 6.35874
R10987 VSS.n889 VSS.n868 6.35874
R10988 VSS.n887 VSS.n870 6.35874
R10989 VSS.n883 VSS.n872 6.35874
R10990 VSS.n890 VSS.n867 6.35874
R10991 VSS.n841 VSS.n789 6.35874
R10992 VSS.n828 VSS.n795 6.35874
R10993 VSS.n827 VSS.n796 6.35874
R10994 VSS.n840 VSS.n790 6.35874
R10995 VSS.n2011 VSS.n1996 6.35874
R10996 VSS.n2016 VSS.n756 6.35874
R10997 VSS.n745 VSS.n721 6.35874
R10998 VSS.n741 VSS.n723 6.35874
R10999 VSS.n737 VSS.n725 6.35874
R11000 VSS.n1359 VSS.n1330 6.35874
R11001 VSS.n679 VSS.n653 6.35874
R11002 VSS.n678 VSS.n654 6.35874
R11003 VSS.n1491 VSS.n1452 6.35874
R11004 VSS.n2163 VSS.n415 6.35874
R11005 VSS.n557 VSS.n554 6.35874
R11006 VSS.n2172 VSS.n409 6.35874
R11007 VSS.n1477 VSS.n1460 6.35874
R11008 VSS.n1485 VSS.n1455 6.35874
R11009 VSS.n440 VSS.n437 6.35874
R11010 VSS.n404 VSS.n403 6.35874
R11011 VSS.n1524 VSS.n1517 6.35874
R11012 VSS.n1537 VSS.n1510 6.35874
R11013 VSS.n2107 VSS.n615 6.35874
R11014 VSS.n2109 VSS.n613 6.35874
R11015 VSS.n2123 VSS.n2120 6.35874
R11016 VSS.n2146 VSS.n607 6.35874
R11017 VSS.n2143 VSS.n2128 6.35874
R11018 VSS.n2140 VSS.n2129 6.35874
R11019 VSS.n2089 VSS.n628 6.35874
R11020 VSS.n2032 VSS.n714 6.3555
R11021 VSS.n2028 VSS.n716 6.3555
R11022 VSS.n695 VSS.n646 6.3555
R11023 VSS.n691 VSS.n647 6.3555
R11024 VSS.n862 VSS.t424 6.32611
R11025 VSS.n2483 VSS.n2477 6.31687
R11026 VSS.n2480 VSS.n2478 6.31687
R11027 VSS.n117 VSS.n112 6.31687
R11028 VSS.n116 VSS.n113 6.31687
R11029 VSS.n146 VSS.n141 6.31687
R11030 VSS.n145 VSS.n142 6.31687
R11031 VSS.n175 VSS.n170 6.31687
R11032 VSS.n174 VSS.n171 6.31687
R11033 VSS.n204 VSS.n199 6.31687
R11034 VSS.n203 VSS.n200 6.31687
R11035 VSS.n233 VSS.n228 6.31687
R11036 VSS.n232 VSS.n229 6.31687
R11037 VSS.n288 VSS.n264 6.31687
R11038 VSS.n287 VSS.n265 6.31687
R11039 VSS.n324 VSS.n319 6.31687
R11040 VSS.n323 VSS.n320 6.31687
R11041 VSS.n3 VSS.n2 6.3142
R11042 VSS.n115 VSS.n114 6.3142
R11043 VSS.n144 VSS.n143 6.3142
R11044 VSS.n173 VSS.n172 6.3142
R11045 VSS.n202 VSS.n201 6.3142
R11046 VSS.n231 VSS.n230 6.3142
R11047 VSS.n286 VSS.n285 6.3142
R11048 VSS.n322 VSS.n321 6.3142
R11049 VSS.n2485 VSS.n2476 6.31016
R11050 VSS.n118 VSS.n111 6.31016
R11051 VSS.n147 VSS.n140 6.31016
R11052 VSS.n176 VSS.n169 6.31016
R11053 VSS.n205 VSS.n198 6.31016
R11054 VSS.n234 VSS.n227 6.31016
R11055 VSS.n289 VSS.n263 6.31016
R11056 VSS.n325 VSS.n318 6.31016
R11057 VSS.n2495 VSS.t64 6.18319
R11058 VSS.n2550 VSS.t338 6.18319
R11059 VSS.n2517 VSS.n2516 6.14978
R11060 VSS.n258 VSS.n257 5.91563
R11061 VSS.n298 VSS.n256 5.91563
R11062 VSS.n28 VSS.n27 5.91466
R11063 VSS.n25 VSS.n24 5.91466
R11064 VSS.n2501 VSS.n2500 5.91466
R11065 VSS.n2504 VSS.n2503 5.91466
R11066 VSS.n294 VSS.n261 5.91289
R11067 VSS.n293 VSS.n292 5.91208
R11068 VSS.n295 VSS.n260 5.91208
R11069 VSS.n468 VSS.t2384 5.79141
R11070 VSS.n498 VSS.t3524 5.79141
R11071 VSS.n485 VSS.t1547 5.79141
R11072 VSS.n83 VSS.t2944 5.79141
R11073 VSS.n1719 VSS.t3790 5.79141
R11074 VSS.n1018 VSS.t2656 5.79141
R11075 VSS.n985 VSS.t4058 5.79141
R11076 VSS.n908 VSS.t3588 5.79141
R11077 VSS.n1853 VSS.t2473 5.79141
R11078 VSS.n898 VSS.t3687 5.79141
R11079 VSS.n853 VSS.t1532 5.79141
R11080 VSS.n861 VSS.t4349 5.79141
R11081 VSS.n863 VSS.t3867 5.79141
R11082 VSS.n793 VSS.t3719 5.79141
R11083 VSS.n799 VSS.t1484 5.79141
R11084 VSS.n785 VSS.t1951 5.79141
R11085 VSS.n757 VSS.t3382 5.79141
R11086 VSS.n2000 VSS.t4099 5.79141
R11087 VSS.n728 VSS.t2134 5.79141
R11088 VSS.n649 VSS.t1329 5.79141
R11089 VSS.n650 VSS.t2267 5.79141
R11090 VSS.n639 VSS.t2949 5.79141
R11091 VSS.n637 VSS.t3315 5.79141
R11092 VSS.n1456 VSS.t3298 5.79141
R11093 VSS.n551 VSS.t1981 5.79141
R11094 VSS.n1454 VSS.t1384 5.79141
R11095 VSS.n398 VSS.t2846 5.79141
R11096 VSS.n627 VSS.t3159 5.79141
R11097 VSS.n625 VSS.t2523 5.79141
R11098 VSS.n621 VSS.t3111 5.79141
R11099 VSS.n619 VSS.t3197 5.79141
R11100 VSS.n611 VSS.t1148 5.79141
R11101 VSS.n2131 VSS.t3909 5.79141
R11102 VSS.n2132 VSS.t4080 5.79141
R11103 VSS.n923 VSS.t2306 5.66271
R11104 VSS.n907 VSS.t3622 5.66271
R11105 VSS.n866 VSS.t2471 5.66271
R11106 VSS.n718 VSS.t3919 5.66271
R11107 VSS.n2130 VSS.t2863 5.66271
R11108 VSS.n541 VSS.n540 5.63259
R11109 VSS.n48 VSS.n47 5.59517
R11110 VSS.n2531 VSS.n2530 5.5328
R11111 VSS.n2421 VSS.n2420 5.52326
R11112 VSS.n532 VSS.n527 5.32359
R11113 VSS.n526 VSS.n525 5.32359
R11114 VSS.n515 VSS.n505 5.32359
R11115 VSS.n504 VSS.n503 5.32359
R11116 VSS.n489 VSS.n486 5.32359
R11117 VSS.n2206 VSS.n379 5.32359
R11118 VSS.n2215 VSS.n372 5.32359
R11119 VSS.t2584 VSS.n2381 5.32359
R11120 VSS.n2290 VSS.t3267 5.32359
R11121 VSS.t3933 VSS.n2281 5.32359
R11122 VSS.n1055 VSS.n1023 5.32359
R11123 VSS.n1092 VSS.t4044 5.32359
R11124 VSS.n1129 VSS.t2334 5.32359
R11125 VSS.n1716 VSS.n1715 5.32359
R11126 VSS.n1678 VSS.t3728 5.32359
R11127 VSS.n1640 VSS.t3959 5.32359
R11128 VSS.n1745 VSS.n980 5.32359
R11129 VSS.n1568 VSS.t2120 5.32359
R11130 VSS.n1605 VSS.t2402 5.32359
R11131 VSS.n952 VSS.n921 5.32359
R11132 VSS.n1777 VSS.n912 5.32359
R11133 VSS.n1162 VSS.t3843 5.32359
R11134 VSS.n1851 VSS.n1850 5.32359
R11135 VSS.n1824 VSS.t3287 5.32359
R11136 VSS.n1192 VSS.t3253 5.32359
R11137 VSS.n1890 VSS.n865 5.32359
R11138 VSS.n1215 VSS.t2355 5.32359
R11139 VSS.n1252 VSS.t2444 5.32359
R11140 VSS.n832 VSS.n794 5.32359
R11141 VSS.n1920 VSS.n781 5.32359
R11142 VSS.n1282 VSS.t1019 5.32359
R11143 VSS.n1994 VSS.n1993 5.32359
R11144 VSS.n1965 VSS.n774 5.32359
R11145 VSS.n1312 VSS.t3080 5.32359
R11146 VSS.n1349 VSS.n1333 5.32359
R11147 VSS.n2030 VSS.n715 5.32359
R11148 VSS.n1383 VSS.t2191 5.32359
R11149 VSS.n2060 VSS.n636 5.32359
R11150 VSS.n688 VSS.n648 5.32359
R11151 VSS.n1413 VSS.t3179 5.32359
R11152 VSS.n2158 VSS.n419 5.32359
R11153 VSS.n1472 VSS.n1464 5.32359
R11154 VSS.n1492 VSS.n1451 5.32359
R11155 VSS.n458 VSS.n457 5.32359
R11156 VSS.n2182 VSS.n399 5.32359
R11157 VSS.n1527 VSS.n1516 5.32359
R11158 VSS.n2125 VSS.n2124 5.32359
R11159 VSS.n2095 VSS.n622 5.32359
R11160 VSS.n1441 VSS.n1430 5.32359
R11161 VSS.n2217 VSS.n2216 5.32359
R11162 VSS.n2249 VSS.n2232 5.32226
R11163 VSS.n2248 VSS.n2233 5.32226
R11164 VSS.n2239 VSS.n2234 5.32226
R11165 VSS.n2318 VSS.n90 5.32226
R11166 VSS.n2330 VSS.n2329 5.32226
R11167 VSS.n2342 VSS.n2331 5.32226
R11168 VSS.n2333 VSS.n2332 5.32226
R11169 VSS.n2412 VSS.n82 5.32226
R11170 VSS.n2391 VSS.t4095 5.32226
R11171 VSS.n2359 VSS.t4277 5.32226
R11172 VSS.n2308 VSS.t2227 5.32226
R11173 VSS.n1046 VSS.t3629 5.32226
R11174 VSS.n1073 VSS.t4024 5.32226
R11175 VSS.n1110 VSS.t1550 5.32226
R11176 VSS.n1730 VSS.n1717 5.32226
R11177 VSS.n1697 VSS.t1242 5.32226
R11178 VSS.n1660 VSS.t4336 5.32226
R11179 VSS.n1007 VSS.n984 5.32226
R11180 VSS.n1759 VSS.n972 5.32226
R11181 VSS.n1586 VSS.t2829 5.32226
R11182 VSS.n941 VSS.n927 5.32226
R11183 VSS.n963 VSS.n915 5.32226
R11184 VSS.n1795 VSS.t967 5.32226
R11185 VSS.n1874 VSS.n1852 5.32226
R11186 VSS.n1838 VSS.n905 5.32226
R11187 VSS.n1806 VSS.t2955 5.32226
R11188 VSS.n885 VSS.n871 5.32226
R11189 VSS.n1902 VSS.n856 5.32226
R11190 VSS.n1233 VSS.t1423 5.32226
R11191 VSS.n823 VSS.n800 5.32226
R11192 VSS.n843 VSS.n788 5.32226
R11193 VSS.n1938 VSS.t1425 5.32226
R11194 VSS.n2012 VSS.n1995 5.32226
R11195 VSS.n1980 VSS.n764 5.32226
R11196 VSS.n1949 VSS.t4255 5.32226
R11197 VSS.n2042 VSS.n708 5.32226
R11198 VSS.n1365 VSS.n1329 5.32226
R11199 VSS.n739 VSS.n724 5.32226
R11200 VSS.n700 VSS.n644 5.32226
R11201 VSS.n2073 VSS.t2653 5.32226
R11202 VSS.n677 VSS.n655 5.32226
R11203 VSS.n561 VSS.n552 5.32226
R11204 VSS.n2168 VSS.n412 5.32226
R11205 VSS.n1480 VSS.n1458 5.32226
R11206 VSS.n442 VSS.n436 5.32226
R11207 VSS.n2195 VSS.n390 5.32226
R11208 VSS.n592 VSS.n459 5.32226
R11209 VSS.n2084 VSS.n631 5.32226
R11210 VSS.n2108 VSS.n614 5.32226
R11211 VSS.n2145 VSS.n2126 5.32226
R11212 VSS.n900 VSS.t3829 5.06876
R11213 VSS.n2522 VSS.n2521 5.0621
R11214 VSS.n2251 VSS.n2250 4.9415
R11215 VSS.n2314 VSS.n2313 4.9415
R11216 VSS.n2349 VSS.n2348 4.9415
R11217 VSS.n2406 VSS.n2405 4.9415
R11218 VSS.n601 VSS.n423 4.9415
R11219 VSS.n2176 VSS.n405 4.9415
R11220 VSS.n2200 VSS.n2199 4.9415
R11221 VSS.n1550 VSS.n373 4.9415
R11222 VSS.n2532 VSS.n2531 4.70661
R11223 VSS.n2493 VSS.n48 4.70569
R11224 VSS.n2463 VSS.n2462 4.61975
R11225 VSS.n106 VSS.n102 4.61975
R11226 VSS.n110 VSS.n109 4.61975
R11227 VSS.n135 VSS.n131 4.61975
R11228 VSS.n139 VSS.n138 4.61975
R11229 VSS.n164 VSS.n160 4.61975
R11230 VSS.n168 VSS.n167 4.61975
R11231 VSS.n193 VSS.n189 4.61975
R11232 VSS.n197 VSS.n196 4.61975
R11233 VSS.n222 VSS.n218 4.61975
R11234 VSS.n226 VSS.n225 4.61975
R11235 VSS.n251 VSS.n247 4.61975
R11236 VSS.n255 VSS.n254 4.61975
R11237 VSS.n313 VSS.n309 4.61975
R11238 VSS.n317 VSS.n316 4.61975
R11239 VSS.n2459 VSS.n55 4.61975
R11240 VSS.t2295 VSS.t1686 4.61698
R11241 VSS.t2488 VSS.t2207 4.61698
R11242 VSS.n2496 VSS.n2495 4.56434
R11243 VSS.n468 VSS.t3846 4.5505
R11244 VSS.n528 VSS.t951 4.5505
R11245 VSS.n528 VSS.t1796 4.5505
R11246 VSS.n498 VSS.t1691 4.5505
R11247 VSS.n485 VSS.t2011 4.5505
R11248 VSS.n83 VSS.t3467 4.5505
R11249 VSS.n1016 VSS.t2516 4.5505
R11250 VSS.n1016 VSS.t3591 4.5505
R11251 VSS.n1719 VSS.t2514 4.5505
R11252 VSS.n1018 VSS.t2170 4.5505
R11253 VSS.n973 VSS.t3203 4.5505
R11254 VSS.n973 VSS.t1656 4.5505
R11255 VSS.n979 VSS.t2743 4.5505
R11256 VSS.n985 VSS.t1308 4.5505
R11257 VSS.n983 VSS.t2891 4.5505
R11258 VSS.n916 VSS.t2397 4.5505
R11259 VSS.n916 VSS.t934 4.5505
R11260 VSS.n924 VSS.t2128 4.5505
R11261 VSS.n928 VSS.t1945 4.5505
R11262 VSS.n928 VSS.t2642 4.5505
R11263 VSS.n929 VSS.t1647 4.5505
R11264 VSS.n926 VSS.t1230 4.5505
R11265 VSS.n926 VSS.t1188 4.5505
R11266 VSS.n925 VSS.t1268 4.5505
R11267 VSS.n925 VSS.t4318 4.5505
R11268 VSS.n919 VSS.t1712 4.5505
R11269 VSS.n908 VSS.t1520 4.5505
R11270 VSS.n903 VSS.t4088 4.5505
R11271 VSS.n896 VSS.t2022 4.5505
R11272 VSS.n896 VSS.t1463 4.5505
R11273 VSS.n1853 VSS.t1335 4.5505
R11274 VSS.n1854 VSS.t3767 4.5505
R11275 VSS.n898 VSS.t2151 4.5505
R11276 VSS.n897 VSS.t3260 4.5505
R11277 VSS.n897 VSS.t4304 4.5505
R11278 VSS.n904 VSS.t3778 4.5505
R11279 VSS.n904 VSS.t2162 4.5505
R11280 VSS.n906 VSS.t2923 4.5505
R11281 VSS.n906 VSS.t3271 4.5505
R11282 VSS.n853 VSS.t1876 4.5505
R11283 VSS.n858 VSS.t2905 4.5505
R11284 VSS.n858 VSS.t2714 4.5505
R11285 VSS.n861 VSS.t2650 4.5505
R11286 VSS.n863 VSS.t4286 4.5505
R11287 VSS.n868 VSS.t3213 4.5505
R11288 VSS.n868 VSS.t3541 4.5505
R11289 VSS.n870 VSS.t2311 4.5505
R11290 VSS.n870 VSS.t1040 4.5505
R11291 VSS.n872 VSS.t2062 4.5505
R11292 VSS.n872 VSS.t3942 4.5505
R11293 VSS.n873 VSS.t1036 4.5505
R11294 VSS.n867 VSS.t2172 4.5505
R11295 VSS.n867 VSS.t1817 4.5505
R11296 VSS.n854 VSS.t1581 4.5505
R11297 VSS.n789 VSS.t2603 4.5505
R11298 VSS.n789 VSS.t1631 4.5505
R11299 VSS.n793 VSS.t984 4.5505
R11300 VSS.n795 VSS.t1380 4.5505
R11301 VSS.n795 VSS.t2946 4.5505
R11302 VSS.n802 VSS.t1059 4.5505
R11303 VSS.n799 VSS.t2362 4.5505
R11304 VSS.n796 VSS.t2190 4.5505
R11305 VSS.n796 VSS.t1015 4.5505
R11306 VSS.n790 VSS.t2222 4.5505
R11307 VSS.n790 VSS.t2115 4.5505
R11308 VSS.n785 VSS.t1861 4.5505
R11309 VSS.n759 VSS.t4041 4.5505
R11310 VSS.n757 VSS.t1275 4.5505
R11311 VSS.n1996 VSS.t2091 4.5505
R11312 VSS.n1996 VSS.t2629 4.5505
R11313 VSS.n2000 VSS.t3329 4.5505
R11314 VSS.n1997 VSS.t3282 4.5505
R11315 VSS.n756 VSS.t1161 4.5505
R11316 VSS.n756 VSS.t4117 4.5505
R11317 VSS.n762 VSS.t4248 4.5505
R11318 VSS.n721 VSS.t1453 4.5505
R11319 VSS.n721 VSS.t1960 4.5505
R11320 VSS.n723 VSS.t3840 4.5505
R11321 VSS.n723 VSS.t3837 4.5505
R11322 VSS.n728 VSS.t2659 4.5505
R11323 VSS.n726 VSS.t3031 4.5505
R11324 VSS.n1330 VSS.t904 4.5505
R11325 VSS.n1330 VSS.t1192 4.5505
R11326 VSS.n638 VSS.t1199 4.5505
R11327 VSS.n649 VSS.t3859 4.5505
R11328 VSS.n653 VSS.t3569 4.5505
R11329 VSS.n653 VSS.t1209 4.5505
R11330 VSS.n656 VSS.t1937 4.5505
R11331 VSS.n654 VSS.t1391 4.5505
R11332 VSS.n654 VSS.t2321 4.5505
R11333 VSS.n650 VSS.t3331 4.5505
R11334 VSS.n645 VSS.t1593 4.5505
R11335 VSS.n639 VSS.t1206 4.5505
R11336 VSS.n637 VSS.t353 4.5505
R11337 VSS.n1452 VSS.t3070 4.5505
R11338 VSS.n1452 VSS.t1316 4.5505
R11339 VSS.n1456 VSS.t1798 4.5505
R11340 VSS.n1463 VSS.t1901 4.5505
R11341 VSS.n415 VSS.t1504 4.5505
R11342 VSS.n415 VSS.t3347 4.5505
R11343 VSS.n553 VSS.t3429 4.5505
R11344 VSS.n551 VSS.t45 4.5505
R11345 VSS.n550 VSS.t3634 4.5505
R11346 VSS.n554 VSS.t3277 4.5505
R11347 VSS.n554 VSS.t127 4.5505
R11348 VSS.n414 VSS.t3097 4.5505
R11349 VSS.n409 VSS.t1404 4.5505
R11350 VSS.n409 VSS.t2610 4.5505
R11351 VSS.n1460 VSS.t1687 4.5505
R11352 VSS.n1460 VSS.t2208 4.5505
R11353 VSS.n1455 VSS.t3052 4.5505
R11354 VSS.n1455 VSS.t1801 4.5505
R11355 VSS.n1454 VSS.t2844 4.5505
R11356 VSS.n1518 VSS.t3501 4.5505
R11357 VSS.n398 VSS.t3054 4.5505
R11358 VSS.n438 VSS.t3733 4.5505
R11359 VSS.n434 VSS.t3691 4.5505
R11360 VSS.n424 VSS.t3517 4.5505
R11361 VSS.n461 VSS.t1972 4.5505
R11362 VSS.n461 VSS.t2981 4.5505
R11363 VSS.n437 VSS.t2271 4.5505
R11364 VSS.n437 VSS.t3129 4.5505
R11365 VSS.n403 VSS.t3531 4.5505
R11366 VSS.n403 VSS.t1622 4.5505
R11367 VSS.n396 VSS.t3370 4.5505
R11368 VSS.n1517 VSS.t2255 4.5505
R11369 VSS.n1517 VSS.t2187 4.5505
R11370 VSS.n1510 VSS.t2842 4.5505
R11371 VSS.n1510 VSS.t2710 4.5505
R11372 VSS.n627 VSS.t2497 4.5505
R11373 VSS.n625 VSS.t4236 4.5505
R11374 VSS.n621 VSS.t1573 4.5505
R11375 VSS.n619 VSS.t3693 4.5505
R11376 VSS.n615 VSS.t2028 4.5505
R11377 VSS.n615 VSS.t656 4.5505
R11378 VSS.n611 VSS.t1575 4.5505
R11379 VSS.n2120 VSS.t3863 4.5505
R11380 VSS.n2120 VSS.t3848 4.5505
R11381 VSS.n607 VSS.t1998 4.5505
R11382 VSS.n607 VSS.t2501 4.5505
R11383 VSS.n2128 VSS.t3007 4.5505
R11384 VSS.n2128 VSS.t4293 4.5505
R11385 VSS.n2129 VSS.t2281 4.5505
R11386 VSS.n2129 VSS.t2030 4.5505
R11387 VSS.n2131 VSS.t1154 4.5505
R11388 VSS.n2132 VSS.t1313 4.5505
R11389 VSS.n606 VSS.t3721 4.5505
R11390 VSS.n606 VSS.t4296 4.5505
R11391 VSS.n618 VSS.t3701 4.5505
R11392 VSS.n628 VSS.t3546 4.5505
R11393 VSS.n628 VSS.t2840 4.5505
R11394 VSS.n109 VSS.n108 4.5005
R11395 VSS.n107 VSS.n106 4.5005
R11396 VSS.n138 VSS.n137 4.5005
R11397 VSS.n136 VSS.n135 4.5005
R11398 VSS.n167 VSS.n166 4.5005
R11399 VSS.n165 VSS.n164 4.5005
R11400 VSS.n196 VSS.n195 4.5005
R11401 VSS.n194 VSS.n193 4.5005
R11402 VSS.n225 VSS.n224 4.5005
R11403 VSS.n223 VSS.n222 4.5005
R11404 VSS.n296 VSS.n295 4.5005
R11405 VSS.n294 VSS.n259 4.5005
R11406 VSS.n293 VSS.n262 4.5005
R11407 VSS.n254 VSS.n253 4.5005
R11408 VSS.n252 VSS.n251 4.5005
R11409 VSS.n316 VSS.n315 4.5005
R11410 VSS.n314 VSS.n313 4.5005
R11411 VSS.n2252 VSS.n2251 4.5005
R11412 VSS.n1145 VSS.n96 4.5005
R11413 VSS.n1624 VSS.n1623 4.5005
R11414 VSS.n1622 VSS.n1621 4.5005
R11415 VSS.n1178 VSS.n1148 4.5005
R11416 VSS.n1542 VSS.n1208 4.5005
R11417 VSS.n1543 VSS.n1268 4.5005
R11418 VSS.n1544 VSS.n1298 4.5005
R11419 VSS.n1545 VSS.n1328 4.5005
R11420 VSS.n1546 VSS.n1399 4.5005
R11421 VSS.n1547 VSS.n1429 4.5005
R11422 VSS.n2078 VSS.n2077 4.5005
R11423 VSS.n1369 VSS.n634 4.5005
R11424 VSS.n1945 VSS.n1944 4.5005
R11425 VSS.n1943 VSS.n1942 4.5005
R11426 VSS.n1237 VSS.n779 4.5005
R11427 VSS.n1802 VSS.n1801 4.5005
R11428 VSS.n1800 VSS.n1799 4.5005
R11429 VSS.n1590 VSS.n910 4.5005
R11430 VSS.n1656 VSS.n1655 4.5005
R11431 VSS.n1114 VSS.n92 4.5005
R11432 VSS.n2313 VSS.n2312 4.5005
R11433 VSS.n1483 VSS.n386 4.5005
R11434 VSS.n1549 VSS.n1508 4.5005
R11435 VSS.n2175 VSS.n2174 4.5005
R11436 VSS.n2052 VSS.n2051 4.5005
R11437 VSS.n2050 VSS.n2049 4.5005
R11438 VSS.n1972 VSS.n704 4.5005
R11439 VSS.n1911 VSS.n1910 4.5005
R11440 VSS.n1909 VSS.n1908 4.5005
R11441 VSS.n1832 VSS.n851 4.5005
R11442 VSS.n1767 VSS.n1766 4.5005
R11443 VSS.n1765 VSS.n1764 4.5005
R11444 VSS.n1688 VSS.n970 4.5005
R11445 VSS.n1082 VSS.n88 4.5005
R11446 VSS.n2350 VSS.n2349 4.5005
R11447 VSS.n2177 VSS.n2176 4.5005
R11448 VSS.n2199 VSS.n2198 4.5005
R11449 VSS.n1551 VSS.n1550 4.5005
R11450 VSS.n601 VSS.n600 4.5005
R11451 VSS.n2155 VSS.n2154 4.5005
R11452 VSS.n684 VSS.n602 4.5005
R11453 VSS.n2025 VSS.n2024 4.5005
R11454 VSS.n2023 VSS.n2022 4.5005
R11455 VSS.n829 VSS.n749 4.5005
R11456 VSS.n1886 VSS.n1885 4.5005
R11457 VSS.n1884 VSS.n1883 4.5005
R11458 VSS.n949 VSS.n892 4.5005
R11459 VSS.n1741 VSS.n1740 4.5005
R11460 VSS.n1739 VSS.n1738 4.5005
R11461 VSS.n1052 VSS.n85 4.5005
R11462 VSS.n2405 VSS.n2404 4.5005
R11463 VSS.n2153 VSS.n2152 4.5005
R11464 VSS.n2103 VSS.n406 4.5005
R11465 VSS.n2080 VSS.n2079 4.5005
R11466 VSS.n1548 VSS.n1450 4.5005
R11467 VSS.n2546 VSS.n2545 4.5005
R11468 VSS.n2529 VSS.n2510 4.5005
R11469 VSS.n2544 VSS.n2543 4.5005
R11470 VSS.n2462 VSS.n2461 4.5005
R11471 VSS.n2460 VSS.n2459 4.5005
R11472 VSS.n357 VSS.n356 4.5005
R11473 VSS.n354 VSS.n97 4.5005
R11474 VSS.n352 VSS.n351 4.5005
R11475 VSS.n350 VSS.n349 4.5005
R11476 VSS.n347 VSS.n343 4.5005
R11477 VSS.n54 VSS.n53 4.5005
R11478 VSS.n2466 VSS.n2465 4.5005
R11479 VSS.n2467 VSS.n52 4.5005
R11480 VSS.n2469 VSS.n2468 4.5005
R11481 VSS.n2470 VSS.n51 4.5005
R11482 VSS.n2472 VSS.n2471 4.5005
R11483 VSS.n2473 VSS.n49 4.5005
R11484 VSS.n2490 VSS.n2489 4.5005
R11485 VSS.n2488 VSS.n50 4.5005
R11486 VSS.n2487 VSS.n2486 4.5005
R11487 VSS.n2484 VSS.n2474 4.5005
R11488 VSS.n2482 VSS.n2481 4.5005
R11489 VSS.n2479 VSS.n1 4.5005
R11490 VSS.n2553 VSS.n2552 4.5005
R11491 VSS.n529 VSS.t2145 4.48817
R11492 VSS.n1017 VSS.t1957 4.48817
R11493 VSS.n976 VSS.t2561 4.48817
R11494 VSS.n918 VSS.t4360 4.48817
R11495 VSS.n930 VSS.t1250 4.48817
R11496 VSS.n894 VSS.t3659 4.48817
R11497 VSS.n895 VSS.t2917 4.48817
R11498 VSS.n860 VSS.t2292 4.48817
R11499 VSS.n874 VSS.t2004 4.48817
R11500 VSS.n869 VSS.t1619 4.48817
R11501 VSS.n791 VSS.t4050 4.48817
R11502 VSS.n797 VSS.t1026 4.48817
R11503 VSS.n798 VSS.t3003 4.48817
R11504 VSS.n787 VSS.t3608 4.48817
R11505 VSS.n1998 VSS.t989 4.48817
R11506 VSS.n753 VSS.t2531 4.48817
R11507 VSS.n1331 VSS.t2245 4.48817
R11508 VSS.n651 VSS.t1701 4.48817
R11509 VSS.n652 VSS.t2648 4.48817
R11510 VSS.n1453 VSS.t4222 4.48817
R11511 VSS.n417 VSS.t3400 4.48817
R11512 VSS.n421 VSS.t3195 4.48817
R11513 VSS.n1466 VSS.t1450 4.48817
R11514 VSS.n1462 VSS.t2024 4.48817
R11515 VSS.n1457 VSS.t3636 4.48817
R11516 VSS.n435 VSS.t4314 4.48817
R11517 VSS.n401 VSS.t2179 4.48817
R11518 VSS.n1519 VSS.t1928 4.48817
R11519 VSS.n1513 VSS.t2807 4.48817
R11520 VSS.n617 VSS.t3528 4.48817
R11521 VSS.n609 VSS.t1543 4.48817
R11522 VSS.n605 VSS.t2583 4.48817
R11523 VSS.n626 VSS.t2825 4.48817
R11524 VSS.n900 VSS.t233 4.0955
R11525 VSS.n901 VSS.t4062 4.0955
R11526 VSS.n901 VSS.t689 4.0955
R11527 VSS.n1019 VSS.t788 4.04494
R11528 VSS.n1019 VSS.t772 4.04494
R11529 VSS.n982 VSS.t2037 4.04494
R11530 VSS.n982 VSS.t2681 4.04494
R11531 VSS.n989 VSS.t2107 4.04494
R11532 VSS.n989 VSS.t2689 4.04494
R11533 VSS.n978 VSS.t2812 4.04494
R11534 VSS.n978 VSS.t2809 4.04494
R11535 VSS.n920 VSS.t2675 4.04494
R11536 VSS.n920 VSS.t1571 4.04494
R11537 VSS.n932 VSS.t2218 4.04494
R11538 VSS.n932 VSS.t2683 4.04494
R11539 VSS.n913 VSS.t284 4.04494
R11540 VSS.n913 VSS.t1814 4.04494
R11541 VSS.n899 VSS.t3559 4.04494
R11542 VSS.n899 VSS.t2679 4.04494
R11543 VSS.n1860 VSS.t2273 4.04494
R11544 VSS.n1860 VSS.t2687 4.04494
R11545 VSS.n876 VSS.t3448 4.04494
R11546 VSS.n876 VSS.t2685 4.04494
R11547 VSS.n859 VSS.t1323 4.04494
R11548 VSS.n859 VSS.t288 4.04494
R11549 VSS.n782 VSS.t864 4.04494
R11550 VSS.n782 VSS.t866 4.04494
R11551 VSS.n809 VSS.t4033 4.04494
R11552 VSS.n809 VSS.t2677 4.04494
R11553 VSS.n777 VSS.t1896 4.04494
R11554 VSS.n777 VSS.t1898 4.04494
R11555 VSS.n776 VSS.t1013 4.04494
R11556 VSS.n776 VSS.t2078 4.04494
R11557 VSS.n775 VSS.t2076 4.04494
R11558 VSS.n775 VSS.t2074 4.04494
R11559 VSS.n763 VSS.t290 4.04494
R11560 VSS.n763 VSS.t2045 4.04494
R11561 VSS.n750 VSS.t712 4.04494
R11562 VSS.n750 VSS.t115 4.04494
R11563 VSS.n2001 VSS.t1556 4.04494
R11564 VSS.n2001 VSS.t2673 4.04494
R11565 VSS.n769 VSS.t282 4.04494
R11566 VSS.n769 VSS.t1333 4.04494
R11567 VSS.n1337 VSS.t870 4.04494
R11568 VSS.n1337 VSS.t860 4.04494
R11569 VSS.n729 VSS.t3581 4.04494
R11570 VSS.n729 VSS.t405 4.04494
R11571 VSS.n717 VSS.t750 4.04494
R11572 VSS.n717 VSS.t666 4.04494
R11573 VSS.n710 VSS.t132 4.04494
R11574 VSS.n710 VSS.t130 4.04494
R11575 VSS.n707 VSS.t140 4.04494
R11576 VSS.n707 VSS.t138 4.04494
R11577 VSS.n643 VSS.t3422 4.04494
R11578 VSS.n643 VSS.t286 4.04494
R11579 VSS.n663 VSS.t1804 4.04494
R11580 VSS.n663 VSS.t395 4.04494
R11581 VSS.n640 VSS.t4207 4.04494
R11582 VSS.n640 VSS.t3641 4.04494
R11583 VSS.n1467 VSS.t3064 4.04494
R11584 VSS.n1467 VSS.t4205 4.04494
R11585 VSS.n420 VSS.t393 4.04494
R11586 VSS.n420 VSS.t1526 4.04494
R11587 VSS.n543 VSS.t3437 4.04494
R11588 VSS.n543 VSS.t403 4.04494
R11589 VSS.n418 VSS.t2816 4.04494
R11590 VSS.n418 VSS.t409 4.04494
R11591 VSS.n388 VSS.t1869 4.04494
R11592 VSS.n388 VSS.t4199 4.04494
R11593 VSS.n400 VSS.t4201 4.04494
R11594 VSS.n400 VSS.t1643 4.04494
R11595 VSS.n430 VSS.t2587 4.04494
R11596 VSS.n430 VSS.t407 4.04494
R11597 VSS.n429 VSS.t1418 4.04494
R11598 VSS.n429 VSS.t397 4.04494
R11599 VSS.n465 VSS.t917 4.04494
R11600 VSS.n465 VSS.t401 4.04494
R11601 VSS.n428 VSS.t3011 4.04494
R11602 VSS.n389 VSS.t4203 4.04494
R11603 VSS.n389 VSS.t1010 4.04494
R11604 VSS.n604 VSS.t371 4.04494
R11605 VSS.n604 VSS.t2453 4.04494
R11606 VSS.n2127 VSS.t3915 4.04494
R11607 VSS.n612 VSS.t3108 4.04494
R11608 VSS.n612 VSS.t4209 4.04494
R11609 VSS.n1022 VSS.t1722 3.8098
R11610 VSS.n1022 VSS.t1718 3.8098
R11611 VSS.n1021 VSS.t1728 3.8098
R11612 VSS.n1021 VSS.t1726 3.8098
R11613 VSS.n1020 VSS.t1732 3.8098
R11614 VSS.n1020 VSS.t1724 3.8098
R11615 VSS.n977 VSS.t2374 3.8098
R11616 VSS.n977 VSS.t2370 3.8098
R11617 VSS.n975 VSS.t2366 3.8098
R11618 VSS.n975 VSS.t2364 3.8098
R11619 VSS.n974 VSS.t2368 3.8098
R11620 VSS.n974 VSS.t2376 3.8098
R11621 VSS.n783 VSS.t298 3.8098
R11622 VSS.n783 VSS.t302 3.8098
R11623 VSS.n784 VSS.t292 3.8098
R11624 VSS.n784 VSS.t296 3.8098
R11625 VSS.n786 VSS.t294 3.8098
R11626 VSS.n786 VSS.t306 3.8098
R11627 VSS.n752 VSS.t2669 3.8098
R11628 VSS.n752 VSS.t2671 3.8098
R11629 VSS.n754 VSS.t2667 3.8098
R11630 VSS.n754 VSS.t2665 3.8098
R11631 VSS.n755 VSS.t2663 3.8098
R11632 VSS.n755 VSS.t2693 3.8098
R11633 VSS.n1332 VSS.t4165 3.8098
R11634 VSS.n1332 VSS.t4167 3.8098
R11635 VSS.n1334 VSS.t4161 3.8098
R11636 VSS.n1334 VSS.t4159 3.8098
R11637 VSS.n1335 VSS.t4163 3.8098
R11638 VSS.n1335 VSS.t4157 3.8098
R11639 VSS.n722 VSS.t332 3.8098
R11640 VSS.n722 VSS.t369 3.8098
R11641 VSS.n720 VSS.t365 3.8098
R11642 VSS.n720 VSS.t334 3.8098
R11643 VSS.n719 VSS.t399 3.8098
R11644 VSS.n719 VSS.t363 3.8098
R11645 VSS.n713 VSS.t760 3.8098
R11646 VSS.n713 VSS.t756 3.8098
R11647 VSS.n712 VSS.t762 3.8098
R11648 VSS.n712 VSS.t758 3.8098
R11649 VSS.n711 VSS.t707 3.8098
R11650 VSS.n711 VSS.t705 3.8098
R11651 VSS.n705 VSS.t872 3.8098
R11652 VSS.n705 VSS.t886 3.8098
R11653 VSS.n1338 VSS.t876 3.8098
R11654 VSS.n1338 VSS.t884 3.8098
R11655 VSS.n1336 VSS.t878 3.8098
R11656 VSS.n1336 VSS.t882 3.8098
R11657 VSS.n355 VSS.t209 3.79962
R11658 VSS.n126 VSS.t627 3.79962
R11659 VSS.n155 VSS.t90 3.79962
R11660 VSS.n184 VSS.t1369 3.79962
R11661 VSS.n213 VSS.t1845 3.79962
R11662 VSS.n242 VSS.t241 3.79962
R11663 VSS.n304 VSS.t574 3.79962
R11664 VSS.n333 VSS.t740 3.79962
R11665 VSS.n2492 VSS.n2491 3.68769
R11666 VSS.n120 VSS.n34 3.68769
R11667 VSS.n149 VSS.n33 3.68769
R11668 VSS.n178 VSS.n35 3.68769
R11669 VSS.n207 VSS.n32 3.68769
R11670 VSS.n236 VSS.n36 3.68769
R11671 VSS.n291 VSS.n37 3.68769
R11672 VSS.n327 VSS.n31 3.68746
R11673 VSS.n2002 VSS.t4138 3.52308
R11674 VSS.n2002 VSS.t1104 3.52308
R11675 VSS.n608 VSS.t20 3.52308
R11676 VSS.n608 VSS.t853 3.52308
R11677 VSS.n2530 VSS.n12 3.488
R11678 VSS.n709 VSS.t659 3.413
R11679 VSS.n709 VSS.t651 3.413
R11680 VSS.n1712 VSS.t4268 3.37782
R11681 VSS.n773 VSS.t160 3.37782
R11682 VSS.n773 VSS.t162 3.37782
R11683 VSS.n772 VSS.t148 3.37782
R11684 VSS.n772 VSS.t146 3.37782
R11685 VSS.n771 VSS.t150 3.37782
R11686 VSS.n771 VSS.t144 3.37782
R11687 VSS.n770 VSS.t172 3.37782
R11688 VSS.n770 VSS.t168 3.37782
R11689 VSS.n768 VSS.t166 3.37782
R11690 VSS.n768 VSS.t170 3.37782
R11691 VSS.n767 VSS.t154 3.37782
R11692 VSS.n767 VSS.t158 3.37782
R11693 VSS.n766 VSS.t156 3.37782
R11694 VSS.n766 VSS.t152 3.37782
R11695 VSS.n623 VSS.t2873 3.37782
R11696 VSS.n610 VSS.t3600 3.37782
R11697 VSS.n2134 VSS.n2133 3.05571
R11698 VSS.n730 VSS.n67 2.97071
R11699 VSS.n353 VSS.n340 2.90641
R11700 VSS.n342 VSS.n341 2.90641
R11701 VSS.n348 VSS.n344 2.90641
R11702 VSS.n346 VSS.n345 2.90641
R11703 VSS.n125 VSS.n98 2.90641
R11704 VSS.n124 VSS.n99 2.90641
R11705 VSS.n123 VSS.n100 2.90641
R11706 VSS.n122 VSS.n101 2.90641
R11707 VSS.n154 VSS.n127 2.90641
R11708 VSS.n153 VSS.n128 2.90641
R11709 VSS.n152 VSS.n129 2.90641
R11710 VSS.n151 VSS.n130 2.90641
R11711 VSS.n183 VSS.n156 2.90641
R11712 VSS.n182 VSS.n157 2.90641
R11713 VSS.n181 VSS.n158 2.90641
R11714 VSS.n180 VSS.n159 2.90641
R11715 VSS.n212 VSS.n185 2.90641
R11716 VSS.n211 VSS.n186 2.90641
R11717 VSS.n210 VSS.n187 2.90641
R11718 VSS.n209 VSS.n188 2.90641
R11719 VSS.n241 VSS.n214 2.90641
R11720 VSS.n240 VSS.n215 2.90641
R11721 VSS.n239 VSS.n216 2.90641
R11722 VSS.n238 VSS.n217 2.90641
R11723 VSS.n303 VSS.n243 2.90641
R11724 VSS.n302 VSS.n244 2.90641
R11725 VSS.n301 VSS.n245 2.90641
R11726 VSS.n300 VSS.n246 2.90641
R11727 VSS.n332 VSS.n305 2.90641
R11728 VSS.n331 VSS.n306 2.90641
R11729 VSS.n330 VSS.n307 2.90641
R11730 VSS.n329 VSS.n308 2.90641
R11731 VSS.n933 VSS.n72 2.86271
R11732 VSS.n1862 VSS.n71 2.86271
R11733 VSS.n877 VSS.n70 2.86271
R11734 VSS.n810 VSS.n69 2.86271
R11735 VSS.n664 VSS.n66 2.86271
R11736 VSS.n575 VSS.n574 2.86271
R11737 VSS.n580 VSS.n579 2.86271
R11738 VSS.n2382 VSS.n76 2.80271
R11739 VSS.n1029 VSS.n75 2.80271
R11740 VSS.n1720 VSS.n74 2.80271
R11741 VSS.n993 VSS.n73 2.80271
R11742 VSS.n2003 VSS.n68 2.80271
R11743 VSS.n855 VSS.t843 2.72794
R11744 VSS.n855 VSS.t1086 2.72794
R11745 VSS.n792 VSS.t3761 2.72794
R11746 VSS.n792 VSS.t2600 2.72794
R11747 VSS.n413 VSS.t324 2.72794
R11748 VSS.n413 VSS.t1448 2.72794
R11749 VSS.n411 VSS.t1319 2.72794
R11750 VSS.n411 VSS.t326 2.72794
R11751 VSS.n2121 VSS.t3796 2.72794
R11752 VSS.n2121 VSS.t3341 2.72794
R11753 VSS.n1449 VSS.n369 2.66271
R11754 VSS.n2253 VSS.n94 2.66171
R11755 VSS.n1144 VSS.n359 2.66171
R11756 VSS.n1625 VSS.n360 2.66171
R11757 VSS.n1620 VSS.n361 2.66171
R11758 VSS.n1177 VSS.n362 2.66171
R11759 VSS.n1207 VSS.n363 2.66171
R11760 VSS.n1267 VSS.n364 2.66171
R11761 VSS.n1297 VSS.n365 2.66171
R11762 VSS.n1327 VSS.n366 2.66171
R11763 VSS.n1398 VSS.n367 2.66171
R11764 VSS.n1428 VSS.n368 2.66171
R11765 VSS.n1507 VSS.n370 2.66171
R11766 VSS.n1541 VSS.n371 2.66171
R11767 VSS.n2511 VSS.t898 2.50972
R11768 VSS.n2527 VSS.t458 2.50972
R11769 VSS.n2525 VSS.t2093 2.50972
R11770 VSS.n2541 VSS.t1401 2.50972
R11771 VSS.n1552 VSS.n0 2.46718
R11772 VSS.n2522 VSS.t2095 2.45409
R11773 VSS.n0 VSS.t2084 2.43747
R11774 VSS.n297 VSS.n296 2.41087
R11775 VSS.n2547 VSS.t1399 2.38597
R11776 VSS.n2548 VSS.n2547 2.36672
R11777 VSS.n105 VSS.n104 2.33691
R11778 VSS.n134 VSS.n133 2.33691
R11779 VSS.n163 VSS.n162 2.33691
R11780 VSS.n192 VSS.n191 2.33691
R11781 VSS.n221 VSS.n220 2.33691
R11782 VSS.n250 VSS.n249 2.33691
R11783 VSS.n312 VSS.n311 2.33691
R11784 VSS.n2458 VSS.n57 2.33691
R11785 VSS.n57 VSS.n56 2.33309
R11786 VSS.n104 VSS.n103 2.33309
R11787 VSS.n133 VSS.n132 2.33309
R11788 VSS.n162 VSS.n161 2.33309
R11789 VSS.n191 VSS.n190 2.33309
R11790 VSS.n220 VSS.n219 2.33309
R11791 VSS.n249 VSS.n248 2.33309
R11792 VSS.n311 VSS.n310 2.33309
R11793 VSS.n2512 VSS.n2511 2.26997
R11794 VSS.n2527 VSS.n2526 2.26997
R11795 VSS.n2525 VSS.n2524 2.26997
R11796 VSS.n2541 VSS.n2540 2.26997
R11797 VSS.n2523 VSS.n2522 2.24629
R11798 VSS.n56 VSS.t217 2.1605
R11799 VSS.n103 VSS.t635 2.1605
R11800 VSS.n132 VSS.t98 2.1605
R11801 VSS.n161 VSS.t1347 2.1605
R11802 VSS.n190 VSS.t1823 2.1605
R11803 VSS.n219 VSS.t249 2.1605
R11804 VSS.n248 VSS.t588 2.1605
R11805 VSS.n310 VSS.t720 2.1605
R11806 VSS.n105 VSS.n58 2.0805
R11807 VSS.n134 VSS.n59 2.0805
R11808 VSS.n163 VSS.n60 2.0805
R11809 VSS.n192 VSS.n61 2.0805
R11810 VSS.n221 VSS.n62 2.0805
R11811 VSS.n250 VSS.n64 2.0805
R11812 VSS.n312 VSS.n63 2.0805
R11813 VSS.n2458 VSS.n2457 2.0805
R11814 VSS.n620 VSS.t3707 2.01032
R11815 VSS.n620 VSS.t3705 2.01032
R11816 VSS.n469 VSS.t2431 1.99806
R11817 VSS.n469 VSS.t2423 1.99806
R11818 VSS.n470 VSS.t2435 1.99806
R11819 VSS.n470 VSS.t2429 1.99806
R11820 VSS.n471 VSS.t2425 1.99806
R11821 VSS.n471 VSS.t2433 1.99806
R11822 VSS.n472 VSS.t2439 1.99806
R11823 VSS.n472 VSS.t2437 1.99806
R11824 VSS.n473 VSS.t2441 1.99806
R11825 VSS.n473 VSS.t2443 1.99806
R11826 VSS.n474 VSS.t2794 1.99806
R11827 VSS.n474 VSS.t2792 1.99806
R11828 VSS.n475 VSS.t3985 1.99806
R11829 VSS.n475 VSS.t2790 1.99806
R11830 VSS.n476 VSS.t3987 1.99806
R11831 VSS.n476 VSS.t3979 1.99806
R11832 VSS.n477 VSS.t3993 1.99806
R11833 VSS.n477 VSS.t3981 1.99806
R11834 VSS.n478 VSS.t3983 1.99806
R11835 VSS.n478 VSS.t3989 1.99806
R11836 VSS.n479 VSS.t3483 1.99806
R11837 VSS.n506 VSS.t1172 1.99806
R11838 VSS.n506 VSS.t1170 1.99806
R11839 VSS.n507 VSS.t445 1.99806
R11840 VSS.n507 VSS.t1176 1.99806
R11841 VSS.n508 VSS.t447 1.99806
R11842 VSS.n508 VSS.t439 1.99806
R11843 VSS.n509 VSS.t437 1.99806
R11844 VSS.n509 VSS.t441 1.99806
R11845 VSS.n499 VSS.t443 1.99806
R11846 VSS.n499 VSS.t449 1.99806
R11847 VSS.n480 VSS.t1736 1.99806
R11848 VSS.n480 VSS.t1740 1.99806
R11849 VSS.n481 VSS.t1779 1.99806
R11850 VSS.n481 VSS.t1738 1.99806
R11851 VSS.n482 VSS.t1783 1.99806
R11852 VSS.n482 VSS.t1787 1.99806
R11853 VSS.n483 VSS.t1777 1.99806
R11854 VSS.n483 VSS.t1789 1.99806
R11855 VSS.n484 VSS.t1791 1.99806
R11856 VSS.n484 VSS.t1781 1.99806
R11857 VSS.n384 VSS.t3133 1.99806
R11858 VSS.n384 VSS.t3137 1.99806
R11859 VSS.n383 VSS.t1440 1.99806
R11860 VSS.n383 VSS.t3135 1.99806
R11861 VSS.n382 VSS.t1428 1.99806
R11862 VSS.n382 VSS.t1434 1.99806
R11863 VSS.n381 VSS.t1442 1.99806
R11864 VSS.n381 VSS.t1436 1.99806
R11865 VSS.n380 VSS.t1438 1.99806
R11866 VSS.n380 VSS.t1430 1.99806
R11867 VSS.n378 VSS.t2578 1.99806
R11868 VSS.n378 VSS.t2576 1.99806
R11869 VSS.n377 VSS.t270 1.99806
R11870 VSS.n377 VSS.t2572 1.99806
R11871 VSS.n376 VSS.t274 1.99806
R11872 VSS.n376 VSS.t278 1.99806
R11873 VSS.n375 VSS.t280 1.99806
R11874 VSS.n375 VSS.t272 1.99806
R11875 VSS.n374 VSS.t238 1.99806
R11876 VSS.n374 VSS.t276 1.99806
R11877 VSS.n81 VSS.t940 1.99806
R11878 VSS.n81 VSS.t946 1.99806
R11879 VSS.n80 VSS.t944 1.99806
R11880 VSS.n80 VSS.t670 1.99806
R11881 VSS.n79 VSS.t668 1.99806
R11882 VSS.n79 VSS.t697 1.99806
R11883 VSS.n78 VSS.t716 1.99806
R11884 VSS.n78 VSS.t701 1.99806
R11885 VSS.n77 VSS.t672 1.99806
R11886 VSS.n77 VSS.t714 1.99806
R11887 VSS.n1024 VSS.t4312 1.99806
R11888 VSS.n1024 VSS.t4310 1.99806
R11889 VSS.n1025 VSS.t4308 1.99806
R11890 VSS.n1025 VSS.t1043 1.99806
R11891 VSS.n1026 VSS.t1057 1.99806
R11892 VSS.n1026 VSS.t1051 1.99806
R11893 VSS.n1027 VSS.t1049 1.99806
R11894 VSS.n1027 VSS.t1055 1.99806
R11895 VSS.n1028 VSS.t1045 1.99806
R11896 VSS.n1028 VSS.t1047 1.99806
R11897 VSS.n1718 VSS.t1766 1.99806
R11898 VSS.n987 VSS.t3810 1.99806
R11899 VSS.n987 VSS.t3812 1.99806
R11900 VSS.n988 VSS.t3814 1.99806
R11901 VSS.n988 VSS.t1851 1.99806
R11902 VSS.n990 VSS.t1605 1.99806
R11903 VSS.n990 VSS.t1599 1.99806
R11904 VSS.n991 VSS.t1953 1.99806
R11905 VSS.n991 VSS.t1603 1.99806
R11906 VSS.n992 VSS.t2080 1.99806
R11907 VSS.n992 VSS.t1991 1.99806
R11908 VSS.n914 VSS.t3407 1.99806
R11909 VSS.n1855 VSS.t1748 1.99806
R11910 VSS.n1855 VSS.t1754 1.99806
R11911 VSS.n1857 VSS.t1752 1.99806
R11912 VSS.n1857 VSS.t320 1.99806
R11913 VSS.n1858 VSS.t318 1.99806
R11914 VSS.n1858 VSS.t312 1.99806
R11915 VSS.n1859 VSS.t310 1.99806
R11916 VSS.n1859 VSS.t316 1.99806
R11917 VSS.n1861 VSS.t322 1.99806
R11918 VSS.n1861 VSS.t308 1.99806
R11919 VSS.n864 VSS.t2039 1.99806
R11920 VSS.n862 VSS.t1264 1.99806
R11921 VSS.n1209 VSS.t2559 1.99806
R11922 VSS.n801 VSS.t1305 1.99806
R11923 VSS.n803 VSS.t1219 1.99806
R11924 VSS.n803 VSS.t1221 1.99806
R11925 VSS.n804 VSS.t1223 1.99806
R11926 VSS.n804 VSS.t49 1.99806
R11927 VSS.n806 VSS.t427 1.99806
R11928 VSS.n806 VSS.t431 1.99806
R11929 VSS.n807 VSS.t433 1.99806
R11930 VSS.n807 VSS.t429 1.99806
R11931 VSS.n808 VSS.t47 1.99806
R11932 VSS.n808 VSS.t51 1.99806
R11933 VSS.n758 VSS.t1277 1.99806
R11934 VSS.n758 VSS.t1076 1.99806
R11935 VSS.n760 VSS.t3141 1.99806
R11936 VSS.n760 VSS.t1341 1.99806
R11937 VSS.n714 VSS.t1095 1.99806
R11938 VSS.n714 VSS.t1099 1.99806
R11939 VSS.n716 VSS.t1097 1.99806
R11940 VSS.n716 VSS.t1093 1.99806
R11941 VSS.n725 VSS.t3586 1.99806
R11942 VSS.n725 VSS.t1102 1.99806
R11943 VSS.n646 VSS.t1127 1.99806
R11944 VSS.n646 VSS.t1114 1.99806
R11945 VSS.n647 VSS.t1125 1.99806
R11946 VSS.n647 VSS.t1120 1.99806
R11947 VSS.n657 VSS.t2993 1.99806
R11948 VSS.n657 VSS.t2991 1.99806
R11949 VSS.n658 VSS.t2989 1.99806
R11950 VSS.n658 VSS.t610 1.99806
R11951 VSS.n660 VSS.t612 1.99806
R11952 VSS.n660 VSS.t910 1.99806
R11953 VSS.n661 VSS.t608 1.99806
R11954 VSS.n661 VSS.t908 1.99806
R11955 VSS.n662 VSS.t906 1.99806
R11956 VSS.n662 VSS.t914 1.99806
R11957 VSS.n1459 VSS.t3372 1.99806
R11958 VSS.n1459 VSS.t2015 1.99806
R11959 VSS.n1461 VSS.t2733 1.99806
R11960 VSS.n1461 VSS.t2304 1.99806
R11961 VSS.n408 VSS.t1933 1.99806
R11962 VSS.n408 VSS.t3050 1.99806
R11963 VSS.n410 VSS.t3883 1.99806
R11964 VSS.n410 VSS.t2297 1.99806
R11965 VSS.n549 VSS.t3749 1.99806
R11966 VSS.n549 VSS.t3743 1.99806
R11967 VSS.n548 VSS.t3745 1.99806
R11968 VSS.n548 VSS.t1685 1.99806
R11969 VSS.n546 VSS.t1679 1.99806
R11970 VSS.n546 VSS.t1681 1.99806
R11971 VSS.n545 VSS.t1673 1.99806
R11972 VSS.n545 VSS.t1677 1.99806
R11973 VSS.n544 VSS.t1683 1.99806
R11974 VSS.n544 VSS.t1671 1.99806
R11975 VSS.n1509 VSS.t37 1.99806
R11976 VSS.n1509 VSS.t29 1.99806
R11977 VSS.n1511 VSS.t31 1.99806
R11978 VSS.n1511 VSS.t41 1.99806
R11979 VSS.n1512 VSS.t43 1.99806
R11980 VSS.n1512 VSS.t35 1.99806
R11981 VSS.n1514 VSS.t39 1.99806
R11982 VSS.n1514 VSS.t927 1.99806
R11983 VSS.n1515 VSS.t923 1.99806
R11984 VSS.n1515 VSS.t921 1.99806
R11985 VSS.n391 VSS.t182 1.99806
R11986 VSS.n391 VSS.t186 1.99806
R11987 VSS.n392 VSS.t174 1.99806
R11988 VSS.n392 VSS.t176 1.99806
R11989 VSS.n394 VSS.t180 1.99806
R11990 VSS.n394 VSS.t184 1.99806
R11991 VSS.n395 VSS.t188 1.99806
R11992 VSS.n395 VSS.t4266 1.99806
R11993 VSS.n397 VSS.t4264 1.99806
R11994 VSS.n397 VSS.t4260 1.99806
R11995 VSS.n460 VSS.t3717 1.99806
R11996 VSS.n462 VSS.t3497 1.99806
R11997 VSS.n462 VSS.t3491 1.99806
R11998 VSS.n463 VSS.t3493 1.99806
R11999 VSS.n463 VSS.t644 1.99806
R12000 VSS.n464 VSS.t662 1.99806
R12001 VSS.n464 VSS.t476 1.99806
R12002 VSS.n466 VSS.t664 1.99806
R12003 VSS.n466 VSS.t474 1.99806
R12004 VSS.n467 VSS.t473 1.99806
R12005 VSS.n467 VSS.t660 1.99806
R12006 VSS.n426 VSS.t754 1.99806
R12007 VSS.n426 VSS.t329 1.99806
R12008 VSS.n453 VSS.t3771 1.99806
R12009 VSS.n453 VSS.t1414 1.99806
R12010 VSS.n431 VSS.t1412 1.99806
R12011 VSS.n431 VSS.t3113 1.99806
R12012 VSS.n432 VSS.t4015 1.99806
R12013 VSS.n432 VSS.t1689 1.99806
R12014 VSS.n1431 VSS.t3877 1.99806
R12015 VSS.n1431 VSS.t2345 1.99806
R12016 VSS.n632 VSS.t2013 1.99806
R12017 VSS.n632 VSS.t2300 1.99806
R12018 VSS.n630 VSS.t1744 1.99806
R12019 VSS.n629 VSS.t999 1.99806
R12020 VSS.n624 VSS.t1286 1.99806
R12021 VSS.n613 VSS.t3604 1.99806
R12022 VSS.n613 VSS.t931 1.99806
R12023 VSS VSS.n2553 1.948
R12024 VSS.n358 VSS.n357 1.7719
R12025 VSS.n2546 VSS.n12 1.5215
R12026 VSS.n691 VSS.n690 1.1975
R12027 VSS.t344 VSS.t70 1.15321
R12028 VSS.t346 VSS.t56 1.15321
R12029 VSS.t342 VSS.t68 1.15321
R12030 VSS.t348 VSS.t62 1.15321
R12031 VSS.t350 VSS.t54 1.15321
R12032 VSS.t354 VSS.t66 1.15321
R12033 VSS.t356 VSS.t60 1.15321
R12034 VSS.t340 VSS.t72 1.15321
R12035 VSS.n2544 VSS.n2510 1.09974
R12036 VSS.n2506 VSS.n2505 1.07796
R12037 VSS.n2509 VSS.n22 1.02303
R12038 VSS.n20 VSS.n19 0.991071
R12039 VSS.n334 VSS.n304 0.921832
R12040 VSS.n2528 VSS.n2527 0.9095
R12041 VSS.n2496 VSS.n29 0.899838
R12042 VSS.n2497 VSS.n28 0.898515
R12043 VSS.n2498 VSS.n25 0.898515
R12044 VSS.n2507 VSS.n2501 0.898515
R12045 VSS.n2506 VSS.n2504 0.898515
R12046 VSS.n121 VSS.n120 0.887926
R12047 VSS.n150 VSS.n149 0.887926
R12048 VSS.n179 VSS.n178 0.887926
R12049 VSS.n208 VSS.n207 0.887926
R12050 VSS.n237 VSS.n236 0.887926
R12051 VSS.n328 VSS.n327 0.887926
R12052 VSS.n20 VSS.n18 0.862992
R12053 VSS.n21 VSS.n15 0.862992
R12054 VSS.n45 VSS.n44 0.862992
R12055 VSS.n46 VSS.n41 0.862992
R12056 VSS.n47 VSS.n38 0.862974
R12057 VSS.n825 VSS.n824 0.85325
R12058 VSS.n335 VSS.n334 0.834479
R12059 VSS.n336 VSS.n335 0.834479
R12060 VSS.n337 VSS.n336 0.834479
R12061 VSS.n338 VSS.n337 0.834479
R12062 VSS.n339 VSS.n338 0.834479
R12063 VSS.n1883 VSS.n893 0.8075
R12064 VSS.n530 VSS.n423 0.80225
R12065 VSS.n356 VSS.n339 0.801983
R12066 VSS.n2542 VSS.n2511 0.7925
R12067 VSS.n936 VSS.n935 0.7895
R12068 VSS.n880 VSS.n879 0.7895
R12069 VSS.n1471 VSS.n1470 0.7895
R12070 VSS.n1521 VSS.n387 0.7895
R12071 VSS.n275 VSS.n274 0.772345
R12072 VSS.n531 VSS.n530 0.7625
R12073 VSS.n2408 VSS.n2407 0.7565
R12074 VSS.n1049 VSS.n1048 0.7565
R12075 VSS.n2106 VSS.n2105 0.74375
R12076 VSS.n2010 VSS.n2009 0.7175
R12077 VSS.n1523 VSS.n1522 0.7175
R12078 VSS.n1881 VSS.n1880 0.6785
R12079 VSS.n827 VSS.n826 0.6785
R12080 VSS.n1488 VSS.n1487 0.6725
R12081 VSS.n2521 VSS.n2520 0.660042
R12082 VSS.n2180 VSS.n2179 0.65825
R12083 VSS.n273 VSS.t2765 0.6505
R12084 VSS.n273 VSS.t2756 0.6505
R12085 VSS.n271 VSS.t2753 0.6505
R12086 VSS.n271 VSS.t2761 0.6505
R12087 VSS.n269 VSS.t2758 0.6505
R12088 VSS.n269 VSS.t2763 0.6505
R12089 VSS.n267 VSS.t2764 0.6505
R12090 VSS.n267 VSS.t2769 0.6505
R12091 VSS.n266 VSS.t2767 0.6505
R12092 VSS.n266 VSS.t2760 0.6505
R12093 VSS.n1736 VSS.n1735 0.64775
R12094 VSS.n890 VSS.n889 0.64775
R12095 VSS.n888 VSS.n887 0.64775
R12096 VSS.n733 VSS.n732 0.63875
R12097 VSS.n557 VSS.n556 0.63125
R12098 VSS.n450 VSS.n449 0.6245
R12099 VSS.n1212 VSS.n1211 0.62075
R12100 VSS.n2333 VSS.n84 0.6185
R12101 VSS.n1473 VSS.n1472 0.61625
R12102 VSS.n2545 VSS.n2509 0.615136
R12103 VSS.n1014 VSS.n1013 0.61325
R12104 VSS.n831 VSS.n830 0.6125
R12105 VSS.n2147 VSS.n2146 0.6095
R12106 VSS.n532 VSS.n531 0.59975
R12107 VSS.n1732 VSS.n1731 0.58775
R12108 VSS.n340 VSS.t226 0.5855
R12109 VSS.n340 VSS.t215 0.5855
R12110 VSS.n341 VSS.t205 0.5855
R12111 VSS.n341 VSS.t224 0.5855
R12112 VSS.n344 VSS.t203 0.5855
R12113 VSS.n344 VSS.t219 0.5855
R12114 VSS.n345 VSS.t211 0.5855
R12115 VSS.n345 VSS.t228 0.5855
R12116 VSS.n2476 VSS.t199 0.5855
R12117 VSS.n2476 VSS.t195 0.5855
R12118 VSS.n2477 VSS.t198 0.5855
R12119 VSS.n2477 VSS.t194 0.5855
R12120 VSS.n2478 VSS.t201 0.5855
R12121 VSS.n2478 VSS.t197 0.5855
R12122 VSS.n2 VSS.t193 0.5855
R12123 VSS.n2 VSS.t200 0.5855
R12124 VSS.n98 VSS.t614 0.5855
R12125 VSS.n98 VSS.t633 0.5855
R12126 VSS.n99 VSS.t623 0.5855
R12127 VSS.n99 VSS.t642 0.5855
R12128 VSS.n100 VSS.t621 0.5855
R12129 VSS.n100 VSS.t637 0.5855
R12130 VSS.n101 VSS.t629 0.5855
R12131 VSS.n101 VSS.t616 0.5855
R12132 VSS.n111 VSS.t1979 0.5855
R12133 VSS.n111 VSS.t1975 0.5855
R12134 VSS.n112 VSS.t1978 0.5855
R12135 VSS.n112 VSS.t1926 0.5855
R12136 VSS.n113 VSS.t1923 0.5855
R12137 VSS.n113 VSS.t1977 0.5855
R12138 VSS.n114 VSS.t1925 0.5855
R12139 VSS.n114 VSS.t1922 0.5855
R12140 VSS.n127 VSS.t77 0.5855
R12141 VSS.n127 VSS.t96 0.5855
R12142 VSS.n128 VSS.t86 0.5855
R12143 VSS.n128 VSS.t75 0.5855
R12144 VSS.n129 VSS.t84 0.5855
R12145 VSS.n129 VSS.t100 0.5855
R12146 VSS.n130 VSS.t92 0.5855
R12147 VSS.n130 VSS.t79 0.5855
R12148 VSS.n140 VSS.t410 0.5855
R12149 VSS.n140 VSS.t416 0.5855
R12150 VSS.n141 VSS.t419 0.5855
R12151 VSS.n141 VSS.t415 0.5855
R12152 VSS.n142 VSS.t412 0.5855
R12153 VSS.n142 VSS.t418 0.5855
R12154 VSS.n143 VSS.t414 0.5855
R12155 VSS.n143 VSS.t411 0.5855
R12156 VSS.n156 VSS.t1356 0.5855
R12157 VSS.n156 VSS.t1345 0.5855
R12158 VSS.n157 VSS.t1365 0.5855
R12159 VSS.n157 VSS.t1354 0.5855
R12160 VSS.n158 VSS.t1363 0.5855
R12161 VSS.n158 VSS.t1349 0.5855
R12162 VSS.n159 VSS.t1371 0.5855
R12163 VSS.n159 VSS.t1358 0.5855
R12164 VSS.n169 VSS.t59 0.5855
R12165 VSS.n169 VSS.t71 0.5855
R12166 VSS.n170 VSS.t57 0.5855
R12167 VSS.n170 VSS.t69 0.5855
R12168 VSS.n171 VSS.t63 0.5855
R12169 VSS.n171 VSS.t55 0.5855
R12170 VSS.n172 VSS.t67 0.5855
R12171 VSS.n172 VSS.t61 0.5855
R12172 VSS.n185 VSS.t1832 0.5855
R12173 VSS.n185 VSS.t1821 0.5855
R12174 VSS.n186 VSS.t1841 0.5855
R12175 VSS.n186 VSS.t1830 0.5855
R12176 VSS.n187 VSS.t1839 0.5855
R12177 VSS.n187 VSS.t1825 0.5855
R12178 VSS.n188 VSS.t1847 0.5855
R12179 VSS.n188 VSS.t1834 0.5855
R12180 VSS.n198 VSS.t118 0.5855
R12181 VSS.n198 VSS.t124 0.5855
R12182 VSS.n199 VSS.t117 0.5855
R12183 VSS.n199 VSS.t123 0.5855
R12184 VSS.n200 VSS.t120 0.5855
R12185 VSS.n200 VSS.t116 0.5855
R12186 VSS.n201 VSS.t122 0.5855
R12187 VSS.n201 VSS.t119 0.5855
R12188 VSS.n214 VSS.t258 0.5855
R12189 VSS.n214 VSS.t247 0.5855
R12190 VSS.n215 VSS.t267 0.5855
R12191 VSS.n215 VSS.t256 0.5855
R12192 VSS.n216 VSS.t265 0.5855
R12193 VSS.n216 VSS.t251 0.5855
R12194 VSS.n217 VSS.t243 0.5855
R12195 VSS.n217 VSS.t260 0.5855
R12196 VSS.n227 VSS.t562 0.5855
R12197 VSS.n227 VSS.t558 0.5855
R12198 VSS.n228 VSS.t561 0.5855
R12199 VSS.n228 VSS.t557 0.5855
R12200 VSS.n229 VSS.t564 0.5855
R12201 VSS.n229 VSS.t560 0.5855
R12202 VSS.n230 VSS.t566 0.5855
R12203 VSS.n230 VSS.t563 0.5855
R12204 VSS.n292 VSS.t596 0.5855
R12205 VSS.n292 VSS.t576 0.5855
R12206 VSS.t2755 VSS.n284 0.5855
R12207 VSS.n284 VSS.t2766 0.5855
R12208 VSS.n282 VSS.t2768 0.5855
R12209 VSS.n282 VSS.t2751 0.5855
R12210 VSS.n280 VSS.t2752 0.5855
R12211 VSS.n280 VSS.t2757 0.5855
R12212 VSS.n278 VSS.t2754 0.5855
R12213 VSS.n278 VSS.t2762 0.5855
R12214 VSS.n276 VSS.t2759 0.5855
R12215 VSS.n276 VSS.t2750 0.5855
R12216 VSS.n261 VSS.t572 0.5855
R12217 VSS.n261 VSS.t584 0.5855
R12218 VSS.n260 VSS.t580 0.5855
R12219 VSS.n260 VSS.t590 0.5855
R12220 VSS.n257 VSS.t594 0.5855
R12221 VSS.n257 VSS.t606 0.5855
R12222 VSS.n256 VSS.t600 0.5855
R12223 VSS.n256 VSS.t582 0.5855
R12224 VSS.t2750 VSS.n263 0.5855
R12225 VSS.t2754 VSS.n263 0.5855
R12226 VSS.t2762 VSS.n264 0.5855
R12227 VSS.t2752 VSS.n264 0.5855
R12228 VSS.t2757 VSS.n265 0.5855
R12229 VSS.t2768 VSS.n265 0.5855
R12230 VSS.n285 VSS.t2751 0.5855
R12231 VSS.n285 VSS.t2755 0.5855
R12232 VSS.n243 VSS.t602 0.5855
R12233 VSS.n243 VSS.t568 0.5855
R12234 VSS.n244 VSS.t586 0.5855
R12235 VSS.n244 VSS.t598 0.5855
R12236 VSS.n245 VSS.t570 0.5855
R12237 VSS.n245 VSS.t592 0.5855
R12238 VSS.n246 VSS.t604 0.5855
R12239 VSS.n246 VSS.t578 0.5855
R12240 VSS.n305 VSS.t730 0.5855
R12241 VSS.n305 VSS.t735 0.5855
R12242 VSS.n306 VSS.t718 0.5855
R12243 VSS.n306 VSS.t727 0.5855
R12244 VSS.n307 VSS.t737 0.5855
R12245 VSS.n307 VSS.t723 0.5855
R12246 VSS.n308 VSS.t732 0.5855
R12247 VSS.n308 VSS.t743 0.5855
R12248 VSS.n318 VSS.t107 0.5855
R12249 VSS.n318 VSS.t110 0.5855
R12250 VSS.n319 VSS.t104 0.5855
R12251 VSS.n319 VSS.t109 0.5855
R12252 VSS.n320 VSS.t112 0.5855
R12253 VSS.n320 VSS.t106 0.5855
R12254 VSS.n321 VSS.t108 0.5855
R12255 VSS.n321 VSS.t111 0.5855
R12256 VSS.n17 VSS.t463 0.5855
R12257 VSS.n17 VSS.t453 0.5855
R12258 VSS.n16 VSS.t377 0.5855
R12259 VSS.n16 VSS.t381 0.5855
R12260 VSS.n14 VSS.t454 0.5855
R12261 VSS.n14 VSS.t456 0.5855
R12262 VSS.n13 VSS.t383 0.5855
R12263 VSS.n13 VSS.t387 0.5855
R12264 VSS.n43 VSS.t460 0.5855
R12265 VSS.n43 VSS.t455 0.5855
R12266 VSS.n42 VSS.t391 0.5855
R12267 VSS.n42 VSS.t385 0.5855
R12268 VSS.n40 VSS.t459 0.5855
R12269 VSS.n40 VSS.t461 0.5855
R12270 VSS.n39 VSS.t389 0.5855
R12271 VSS.n39 VSS.t373 0.5855
R12272 VSS.n27 VSS.t889 0.5855
R12273 VSS.n27 VSS.t887 0.5855
R12274 VSS.n26 VSS.t347 0.5855
R12275 VSS.n26 VSS.t343 0.5855
R12276 VSS.n24 VSS.t890 0.5855
R12277 VSS.n24 VSS.t891 0.5855
R12278 VSS.n23 VSS.t349 0.5855
R12279 VSS.n23 VSS.t351 0.5855
R12280 VSS.n2500 VSS.t892 0.5855
R12281 VSS.n2500 VSS.t893 0.5855
R12282 VSS.n2499 VSS.t355 0.5855
R12283 VSS.n2499 VSS.t357 0.5855
R12284 VSS.n2503 VSS.t896 0.5855
R12285 VSS.n2503 VSS.t894 0.5855
R12286 VSS.n2502 VSS.t341 0.5855
R12287 VSS.n2502 VSS.t337 0.5855
R12288 VSS.n735 VSS.n734 0.57875
R12289 VSS.n961 VSS.n960 0.57575
R12290 VSS.n2052 VSS.n703 0.5495
R12291 VSS.n842 VSS.n841 0.54575
R12292 VSS.n1837 VSS.n1836 0.545
R12293 VSS.n682 VSS.n681 0.54125
R12294 VSS.n2093 VSS.n2092 0.5375
R12295 VSS.n2413 VSS.n2412 0.5345
R12296 VSS.n2215 VSS.n2214 0.5345
R12297 VSS.n2065 VSS.n2064 0.52925
R12298 VSS.n835 VSS.n834 0.5285
R12299 VSS.n680 VSS.n679 0.5105
R12300 VSS.n2088 VSS.n2087 0.5105
R12301 VSS.n1744 VSS.n1743 0.5075
R12302 VSS.n2056 VSS.n2055 0.50525
R12303 VSS.n2112 VSS.n2111 0.5045
R12304 VSS.n2094 VSS.n2093 0.4985
R12305 VSS.n959 VSS.n958 0.4955
R12306 VSS.n1474 VSS.n1473 0.4955
R12307 VSS.n445 VSS.n444 0.4955
R12308 VSS.n2161 VSS.n2160 0.49025
R12309 VSS.n446 VSS.n445 0.4775
R12310 VSS.n1981 VSS.n1980 0.47525
R12311 VSS.n2545 VSS.n2544 0.474546
R12312 VSS.n701 VSS.n700 0.4745
R12313 VSS.n1889 VSS.n1888 0.47075
R12314 VSS.n738 VSS.n737 0.46925
R12315 VSS.n599 VSS.n598 0.4685
R12316 VSS.n2163 VSS.n2162 0.46325
R12317 VSS.n1901 VSS.n1900 0.46175
R12318 VSS.n937 VSS.n936 0.45725
R12319 VSS.n881 VSS.n880 0.45725
R12320 VSS.n1484 VSS.n1483 0.4535
R12321 VSS.n1449 VSS.n1448 0.4535
R12322 VSS.n1007 VSS.n1006 0.4505
R12323 VSS.n489 VSS.n488 0.44975
R12324 VSS.n1009 VSS.n1008 0.44675
R12325 VSS.n1984 VSS.n1983 0.44225
R12326 VSS.n1896 VSS.n1895 0.4415
R12327 VSS.n1550 VSS.n1549 0.4415
R12328 VSS.n1549 VSS.n1548 0.4415
R12329 VSS.n1548 VSS.n1547 0.4415
R12330 VSS.n1547 VSS.n1546 0.4415
R12331 VSS.n1546 VSS.n1545 0.4415
R12332 VSS.n1545 VSS.n1544 0.4415
R12333 VSS.n1544 VSS.n1543 0.4415
R12334 VSS.n1543 VSS.n1542 0.4415
R12335 VSS.n1542 VSS.n1148 0.4415
R12336 VSS.n1622 VSS.n1148 0.4415
R12337 VSS.n1623 VSS.n1622 0.4415
R12338 VSS.n1623 VSS.n96 0.4415
R12339 VSS.n2251 VSS.n96 0.4415
R12340 VSS.n2199 VSS.n386 0.4415
R12341 VSS.n2079 VSS.n386 0.4415
R12342 VSS.n2079 VSS.n2078 0.4415
R12343 VSS.n2078 VSS.n634 0.4415
R12344 VSS.n1944 VSS.n634 0.4415
R12345 VSS.n1944 VSS.n1943 0.4415
R12346 VSS.n1943 VSS.n779 0.4415
R12347 VSS.n1801 VSS.n779 0.4415
R12348 VSS.n1801 VSS.n1800 0.4415
R12349 VSS.n1800 VSS.n910 0.4415
R12350 VSS.n1655 VSS.n910 0.4415
R12351 VSS.n1655 VSS.n92 0.4415
R12352 VSS.n2313 VSS.n92 0.4415
R12353 VSS.n2176 VSS.n2175 0.4415
R12354 VSS.n2175 VSS.n406 0.4415
R12355 VSS.n2051 VSS.n406 0.4415
R12356 VSS.n2051 VSS.n2050 0.4415
R12357 VSS.n2050 VSS.n704 0.4415
R12358 VSS.n1910 VSS.n704 0.4415
R12359 VSS.n1910 VSS.n1909 0.4415
R12360 VSS.n1909 VSS.n851 0.4415
R12361 VSS.n1766 VSS.n851 0.4415
R12362 VSS.n1766 VSS.n1765 0.4415
R12363 VSS.n1765 VSS.n970 0.4415
R12364 VSS.n970 VSS.n88 0.4415
R12365 VSS.n2349 VSS.n88 0.4415
R12366 VSS.n2154 VSS.n601 0.4415
R12367 VSS.n2154 VSS.n2153 0.4415
R12368 VSS.n2153 VSS.n602 0.4415
R12369 VSS.n2024 VSS.n602 0.4415
R12370 VSS.n2024 VSS.n2023 0.4415
R12371 VSS.n2023 VSS.n749 0.4415
R12372 VSS.n1885 VSS.n749 0.4415
R12373 VSS.n1885 VSS.n1884 0.4415
R12374 VSS.n1884 VSS.n892 0.4415
R12375 VSS.n1740 VSS.n892 0.4415
R12376 VSS.n1740 VSS.n1739 0.4415
R12377 VSS.n1739 VSS.n85 0.4415
R12378 VSS.n2405 VSS.n85 0.4415
R12379 VSS.n1491 VSS.n1490 0.43925
R12380 VSS.n948 VSS.n947 0.43475
R12381 VSS.n840 VSS.n839 0.43325
R12382 VSS.n2172 VSS.n2171 0.43325
R12383 VSS.n2149 VSS.n2148 0.43325
R12384 VSS.n1476 VSS.n1475 0.43175
R12385 VSS.n2146 VSS.n2145 0.43175
R12386 VSS.n1747 VSS.n1746 0.422
R12387 VSS.n1727 VSS.n1726 0.4205
R12388 VSS.n2008 VSS.n2007 0.4205
R12389 VSS.n2140 VSS.n2139 0.41075
R12390 VSS.n2103 VSS.n2102 0.39725
R12391 VSS.n540 VSS.n539 0.3965
R12392 VSS.n1842 VSS.n1841 0.39425
R12393 VSS.n1988 VSS.n1987 0.39425
R12394 VSS.n591 VSS.n590 0.3935
R12395 VSS.n1480 VSS.n1479 0.3905
R12396 VSS.n2183 VSS.n2182 0.3905
R12397 VSS.n2547 VSS.n2546 0.3875
R12398 VSS.n821 VSS.n820 0.3875
R12399 VSS.n2529 VSS.n2528 0.3875
R12400 VSS.n2543 VSS.n2542 0.3875
R12401 VSS.n2091 VSS.n2090 0.38375
R12402 VSS.n939 VSS.n938 0.3815
R12403 VSS.n938 VSS.n937 0.3815
R12404 VSS.n883 VSS.n882 0.3815
R12405 VSS.n882 VSS.n881 0.3815
R12406 VSS.n947 VSS.n946 0.37925
R12407 VSS.n2090 VSS.n2089 0.37925
R12408 VSS.n951 VSS.n950 0.37625
R12409 VSS.n887 VSS.n886 0.374
R12410 VSS.n1877 VSS.n1876 0.37025
R12411 VSS.n2254 VSS.n2253 0.3695
R12412 VSS.n1144 VSS.n1143 0.3695
R12413 VSS.n1626 VSS.n1625 0.3695
R12414 VSS.n1620 VSS.n1619 0.3695
R12415 VSS.n1177 VSS.n1176 0.3695
R12416 VSS.n1207 VSS.n1206 0.3695
R12417 VSS.n1267 VSS.n1266 0.3695
R12418 VSS.n1297 VSS.n1296 0.3695
R12419 VSS.n1327 VSS.n1326 0.3695
R12420 VSS.n2015 VSS.n2014 0.3695
R12421 VSS.n2007 VSS.n2006 0.3695
R12422 VSS.n1398 VSS.n1397 0.3695
R12423 VSS.n1428 VSS.n1427 0.3695
R12424 VSS.n1507 VSS.n1506 0.3695
R12425 VSS.n517 VSS.n516 0.3695
R12426 VSS.n275 VSS.n262 0.36721
R12427 VSS.n2248 VSS.n2247 0.3665
R12428 VSS.n2239 VSS.n2238 0.3665
R12429 VSS.n2319 VSS.n2318 0.3665
R12430 VSS.n2329 VSS.n2328 0.3665
R12431 VSS.n2342 VSS.n2341 0.3665
R12432 VSS.n2124 VSS.n2119 0.3665
R12433 VSS.n490 VSS.n489 0.3665
R12434 VSS.n503 VSS.n502 0.3665
R12435 VSS.n525 VSS.n524 0.3665
R12436 VSS.n676 VSS.n675 0.365
R12437 VSS.n1751 VSS.n1750 0.3635
R12438 VSS.n1894 VSS.n1893 0.3635
R12439 VSS.n2047 VSS.n2046 0.3635
R12440 VSS.n2037 VSS.n2036 0.3635
R12441 VSS.n2027 VSS.n2026 0.3635
R12442 VSS.n2156 VSS.n2155 0.3605
R12443 VSS.n564 VSS.n563 0.3605
R12444 VSS.n2532 VSS.n2518 0.350882
R12445 VSS.n1904 VSS.n1903 0.35075
R12446 VSS.n2122 VSS.n603 0.35075
R12447 VSS.n944 VSS.n943 0.34925
R12448 VSS.n2164 VSS.n2163 0.34925
R12449 VSS.n2178 VSS.n2177 0.3485
R12450 VSS.n963 VSS.n962 0.34775
R12451 VSS.n1840 VSS.n1839 0.34775
R12452 VSS.n1985 VSS.n1984 0.34775
R12453 VSS.n2012 VSS.n2011 0.34775
R12454 VSS.n694 VSS.n693 0.34775
R12455 VSS.n2108 VSS.n2107 0.34775
R12456 VSS.n299 VSS.n298 0.344331
R12457 VSS.n2521 VSS.n2510 0.344011
R12458 VSS.n687 VSS.n686 0.344
R12459 VSS.n1891 VSS.n1890 0.3395
R12460 VSS.n2031 VSS.n2030 0.3395
R12461 VSS.n1733 VSS.n1732 0.33725
R12462 VSS.n2247 VSS.n2246 0.3365
R12463 VSS.n2246 VSS.n2245 0.3365
R12464 VSS.n2245 VSS.n2244 0.3365
R12465 VSS.n2244 VSS.n2243 0.3365
R12466 VSS.n2243 VSS.n2242 0.3365
R12467 VSS.n2242 VSS.n2241 0.3365
R12468 VSS.n2241 VSS.n2240 0.3365
R12469 VSS.n2238 VSS.n2237 0.3365
R12470 VSS.n2237 VSS.n2236 0.3365
R12471 VSS.n2236 VSS.n2235 0.3365
R12472 VSS.n2235 VSS.n91 0.3365
R12473 VSS.n2316 VSS.n2315 0.3365
R12474 VSS.n2317 VSS.n2316 0.3365
R12475 VSS.n2320 VSS.n2319 0.3365
R12476 VSS.n2321 VSS.n2320 0.3365
R12477 VSS.n2322 VSS.n2321 0.3365
R12478 VSS.n2323 VSS.n2322 0.3365
R12479 VSS.n2324 VSS.n2323 0.3365
R12480 VSS.n2325 VSS.n2324 0.3365
R12481 VSS.n2326 VSS.n2325 0.3365
R12482 VSS.n2328 VSS.n2327 0.3365
R12483 VSS.n2327 VSS.n89 0.3365
R12484 VSS.n2347 VSS.n2346 0.3365
R12485 VSS.n2346 VSS.n2345 0.3365
R12486 VSS.n2345 VSS.n2344 0.3365
R12487 VSS.n2344 VSS.n2343 0.3365
R12488 VSS.n2341 VSS.n2340 0.3365
R12489 VSS.n2340 VSS.n2339 0.3365
R12490 VSS.n2339 VSS.n2338 0.3365
R12491 VSS.n2338 VSS.n2337 0.3365
R12492 VSS.n2337 VSS.n2336 0.3365
R12493 VSS.n2336 VSS.n2335 0.3365
R12494 VSS.n2335 VSS.n2334 0.3365
R12495 VSS.n2409 VSS.n2408 0.3365
R12496 VSS.n2410 VSS.n2409 0.3365
R12497 VSS.n2411 VSS.n2410 0.3365
R12498 VSS.n2415 VSS.n2414 0.3365
R12499 VSS.n2416 VSS.n2415 0.3365
R12500 VSS.n2417 VSS.n2416 0.3365
R12501 VSS.n2418 VSS.n2417 0.3365
R12502 VSS.n2419 VSS.n2418 0.3365
R12503 VSS.n2420 VSS.n2419 0.3365
R12504 VSS.n2390 VSS.n2389 0.3365
R12505 VSS.n2389 VSS.n2388 0.3365
R12506 VSS.n2388 VSS.n2387 0.3365
R12507 VSS.n2387 VSS.n2386 0.3365
R12508 VSS.n2386 VSS.n2385 0.3365
R12509 VSS.n2385 VSS.n2384 0.3365
R12510 VSS.n2384 VSS.n2383 0.3365
R12511 VSS.n2383 VSS.n2382 0.3365
R12512 VSS.n1072 VSS.n1071 0.3365
R12513 VSS.n1054 VSS.n1053 0.3365
R12514 VSS.n1051 VSS.n1050 0.3365
R12515 VSS.n1050 VSS.n1049 0.3365
R12516 VSS.n1048 VSS.n1047 0.3365
R12517 VSS.n1045 VSS.n1044 0.3365
R12518 VSS.n1699 VSS.n1698 0.3365
R12519 VSS.n1711 VSS.n1710 0.3365
R12520 VSS.n1725 VSS.n1724 0.3365
R12521 VSS.n1724 VSS.n1723 0.3365
R12522 VSS.n1723 VSS.n1722 0.3365
R12523 VSS.n1722 VSS.n1721 0.3365
R12524 VSS.n1721 VSS.n1720 0.3365
R12525 VSS.n1567 VSS.n1566 0.3365
R12526 VSS.n1566 VSS.n1565 0.3365
R12527 VSS.n1565 VSS.n1564 0.3365
R12528 VSS.n1564 VSS.n971 0.3365
R12529 VSS.n1763 VSS.n1762 0.3365
R12530 VSS.n1762 VSS.n1761 0.3365
R12531 VSS.n1761 VSS.n1760 0.3365
R12532 VSS.n1755 VSS.n1754 0.3365
R12533 VSS.n1752 VSS.n1751 0.3365
R12534 VSS.n1750 VSS.n1749 0.3365
R12535 VSS.n1004 VSS.n1003 0.3365
R12536 VSS.n997 VSS.n996 0.3365
R12537 VSS.n1794 VSS.n1793 0.3365
R12538 VSS.n968 VSS.n967 0.3365
R12539 VSS.n1829 VSS.n1828 0.3365
R12540 VSS.n1830 VSS.n1829 0.3365
R12541 VSS.n1871 VSS.n1870 0.3365
R12542 VSS.n1868 VSS.n1867 0.3365
R12543 VSS.n1867 VSS.n1866 0.3365
R12544 VSS.n1863 VSS.n1862 0.3365
R12545 VSS.n1214 VSS.n1213 0.3365
R12546 VSS.n1210 VSS.n852 0.3365
R12547 VSS.n1937 VSS.n1936 0.3365
R12548 VSS.n1914 VSS.n1913 0.3365
R12549 VSS.n849 VSS.n848 0.3365
R12550 VSS.n846 VSS.n845 0.3365
R12551 VSS.n818 VSS.n817 0.3365
R12552 VSS.n815 VSS.n814 0.3365
R12553 VSS.n1951 VSS.n1950 0.3365
R12554 VSS.n1958 VSS.n1957 0.3365
R12555 VSS.n1967 VSS.n1966 0.3365
R12556 VSS.n1968 VSS.n1967 0.3365
R12557 VSS.n1969 VSS.n1968 0.3365
R12558 VSS.n1977 VSS.n1976 0.3365
R12559 VSS.n1978 VSS.n1977 0.3365
R12560 VSS.n1987 VSS.n1986 0.3365
R12561 VSS.n2021 VSS.n2020 0.3365
R12562 VSS.n2018 VSS.n2017 0.3365
R12563 VSS.n2004 VSS.n2003 0.3365
R12564 VSS.n1382 VSS.n1381 0.3365
R12565 VSS.n1364 VSS.n1363 0.3365
R12566 VSS.n1358 VSS.n1357 0.3365
R12567 VSS.n1355 VSS.n1354 0.3365
R12568 VSS.n1348 VSS.n1347 0.3365
R12569 VSS.n2046 VSS.n2045 0.3365
R12570 VSS.n2036 VSS.n2035 0.3365
R12571 VSS.n2035 VSS.n2034 0.3365
R12572 VSS.n2034 VSS.n2033 0.3365
R12573 VSS.n747 VSS.n746 0.3365
R12574 VSS.n744 VSS.n743 0.3365
R12575 VSS.n2072 VSS.n2071 0.3365
R12576 VSS.n2063 VSS.n2062 0.3365
R12577 VSS.n672 VSS.n671 0.3365
R12578 VSS.n669 VSS.n668 0.3365
R12579 VSS.n1479 VSS.n1478 0.3365
R12580 VSS.n567 VSS.n566 0.3365
R12581 VSS.n570 VSS.n569 0.3365
R12582 VSS.n1536 VSS.n1535 0.3365
R12583 VSS.n1533 VSS.n1532 0.3365
R12584 VSS.n2193 VSS.n2192 0.3365
R12585 VSS.n2192 VSS.n2191 0.3365
R12586 VSS.n2191 VSS.n2190 0.3365
R12587 VSS.n2190 VSS.n2189 0.3365
R12588 VSS.n588 VSS.n587 0.3365
R12589 VSS.n583 VSS.n582 0.3365
R12590 VSS.n1448 VSS.n1447 0.3365
R12591 VSS.n1447 VSS.n1446 0.3365
R12592 VSS.n1446 VSS.n1445 0.3365
R12593 VSS.n1445 VSS.n1444 0.3365
R12594 VSS.n1444 VSS.n1443 0.3365
R12595 VSS.n1443 VSS.n1442 0.3365
R12596 VSS.n1440 VSS.n1439 0.3365
R12597 VSS.n1439 VSS.n1438 0.3365
R12598 VSS.n1438 VSS.n1437 0.3365
R12599 VSS.n1433 VSS.n1432 0.3365
R12600 VSS.n2115 VSS.n2114 0.3365
R12601 VSS.n2213 VSS.n2212 0.3365
R12602 VSS.n2212 VSS.n2211 0.3365
R12603 VSS.n2211 VSS.n2210 0.3365
R12604 VSS.n2210 VSS.n2209 0.3365
R12605 VSS.n2209 VSS.n2208 0.3365
R12606 VSS.n2208 VSS.n2207 0.3365
R12607 VSS.n2205 VSS.n2204 0.3365
R12608 VSS.n2204 VSS.n2203 0.3365
R12609 VSS.n2203 VSS.n2202 0.3365
R12610 VSS.n2202 VSS.n2201 0.3365
R12611 VSS.n487 VSS.n385 0.3365
R12612 VSS.n491 VSS.n490 0.3365
R12613 VSS.n492 VSS.n491 0.3365
R12614 VSS.n493 VSS.n492 0.3365
R12615 VSS.n494 VSS.n493 0.3365
R12616 VSS.n495 VSS.n494 0.3365
R12617 VSS.n496 VSS.n495 0.3365
R12618 VSS.n497 VSS.n496 0.3365
R12619 VSS.n502 VSS.n501 0.3365
R12620 VSS.n501 VSS.n500 0.3365
R12621 VSS.n511 VSS.n510 0.3365
R12622 VSS.n512 VSS.n511 0.3365
R12623 VSS.n513 VSS.n512 0.3365
R12624 VSS.n514 VSS.n513 0.3365
R12625 VSS.n518 VSS.n517 0.3365
R12626 VSS.n519 VSS.n518 0.3365
R12627 VSS.n520 VSS.n519 0.3365
R12628 VSS.n521 VSS.n520 0.3365
R12629 VSS.n522 VSS.n521 0.3365
R12630 VSS.n523 VSS.n522 0.3365
R12631 VSS.n534 VSS.n533 0.3365
R12632 VSS.n535 VSS.n534 0.3365
R12633 VSS.n536 VSS.n535 0.3365
R12634 VSS.n537 VSS.n536 0.3365
R12635 VSS.n538 VSS.n537 0.3365
R12636 VSS.n539 VSS.n538 0.3365
R12637 VSS.n819 VSS.n818 0.33425
R12638 VSS.n673 VSS.n672 0.33425
R12639 VSS.n566 VSS.n565 0.33425
R12640 VSS.n592 VSS.n591 0.3335
R12641 VSS.n2096 VSS.n2095 0.3335
R12642 VSS.n516 VSS.n515 0.3335
R12643 VSS.n1477 VSS.n1476 0.33125
R12644 VSS.n1756 VSS.n1755 0.32825
R12645 VSS.n1900 VSS.n1899 0.32825
R12646 VSS.n950 VSS.n949 0.3275
R12647 VSS.n524 VSS.n423 0.3275
R12648 VSS.n1844 VSS.n1843 0.32675
R12649 VSS.n746 VSS.n745 0.326
R12650 VSS.n560 VSS.n559 0.32525
R12651 VSS.n2187 VSS.n2186 0.32525
R12652 VSS.n2101 VSS.n2100 0.32525
R12653 VSS.n2145 VSS.n2144 0.32525
R12654 VSS.n2166 VSS.n2165 0.3245
R12655 VSS.n1357 VSS.n1356 0.32375
R12656 VSS.n1490 VSS.n1489 0.32375
R12657 VSS.n440 VSS.n439 0.32
R12658 VSS.n1481 VSS.n1480 0.31925
R12659 VSS.n1839 VSS.n1838 0.31775
R12660 VSS.n561 VSS.n560 0.31775
R12661 VSS.n1525 VSS.n1524 0.31775
R12662 VSS.n442 VSS.n441 0.31775
R12663 VSS.n837 VSS.n836 0.31475
R12664 VSS.n597 VSS.n596 0.314
R12665 VSS.n1726 VSS.n1725 0.3125
R12666 VSS.n2136 VSS.n2135 0.3095
R12667 VSS.n1874 VSS.n1873 0.3065
R12668 VSS.n2159 VSS.n2158 0.3065
R12669 VSS.n593 VSS.n592 0.3065
R12670 VSS.n2109 VSS.n2108 0.3065
R12671 VSS.n2022 VSS.n751 0.3035
R12672 VSS.n2142 VSS.n2141 0.3035
R12673 VSS.n1846 VSS.n1845 0.30275
R12674 VSS.n2162 VSS.n2161 0.29975
R12675 VSS.n2155 VSS.n422 0.29825
R12676 VSS.n277 VSS.n275 0.297779
R12677 VSS.n945 VSS.n944 0.2975
R12678 VSS.n1834 VSS.n1833 0.296
R12679 VSS.n1478 VSS.n1477 0.29375
R12680 VSS.n598 VSS.n597 0.29225
R12681 VSS.n2033 VSS.n2032 0.2915
R12682 VSS.n741 VSS.n740 0.29
R12683 VSS.n1011 VSS.n1010 0.28775
R12684 VSS.n1845 VSS.n1844 0.28625
R12685 VSS.n115 VSS.n10 0.28617
R12686 VSS.n144 VSS.n9 0.28617
R12687 VSS.n173 VSS.n8 0.28617
R12688 VSS.n202 VSS.n7 0.28617
R12689 VSS.n231 VSS.n6 0.28617
R12690 VSS.n286 VSS.n4 0.28617
R12691 VSS.n322 VSS.n5 0.28617
R12692 VSS.n1714 VSS.n1713 0.2855
R12693 VSS.n1729 VSS.n1728 0.2855
R12694 VSS.n1003 VSS.n1002 0.2855
R12695 VSS.n814 VSS.n813 0.2855
R12696 VSS.n668 VSS.n667 0.2855
R12697 VSS.n571 VSS.n570 0.2855
R12698 VSS.n2201 VSS.n2200 0.2855
R12699 VSS.n2177 VSS.n404 0.28325
R12700 VSS.n1055 VSS.n1054 0.2825
R12701 VSS.n1731 VSS.n1730 0.2825
R12702 VSS.n1777 VSS.n1776 0.2825
R12703 VSS.n1920 VSS.n1919 0.2825
R12704 VSS.n2085 VSS.n2084 0.2825
R12705 VSS.n2206 VSS.n2205 0.2825
R12706 VSS.n1008 VSS.n1007 0.28025
R12707 VSS.n1745 VSS.n1744 0.2795
R12708 VSS.n1012 VSS.n1011 0.2795
R12709 VSS.n935 VSS.n934 0.2795
R12710 VSS.n1865 VSS.n1864 0.2795
R12711 VSS.n1899 VSS.n1898 0.2795
R12712 VSS.n879 VSS.n878 0.2795
R12713 VSS.n2006 VSS.n2005 0.2795
R12714 VSS.n2040 VSS.n2039 0.2795
R12715 VSS.n731 VSS.n730 0.2795
R12716 VSS.n2160 VSS.n2159 0.2795
R12717 VSS.n452 VSS.n451 0.2795
R12718 VSS.n2111 VSS.n2110 0.2795
R12719 VSS.n955 VSS.n954 0.27875
R12720 VSS.n1971 VSS.n1970 0.27875
R12721 VSS.n2157 VSS.n2156 0.27875
R12722 VSS.n2181 VSS.n2180 0.27875
R12723 VSS.n1919 VSS.n1918 0.27725
R12724 VSS.n2185 VSS.n2184 0.27725
R12725 VSS.n1041 VSS.n1040 0.2765
R12726 VSS.n1039 VSS.n1038 0.2765
R12727 VSS.n1037 VSS.n1036 0.2765
R12728 VSS.n1035 VSS.n1034 0.2765
R12729 VSS.n1033 VSS.n1032 0.2765
R12730 VSS.n1031 VSS.n1030 0.2765
R12731 VSS.n1738 VSS.n1015 0.2765
R12732 VSS.n995 VSS.n994 0.2765
R12733 VSS.n1468 VSS.n407 0.2765
R12734 VSS.n584 VSS.n583 0.2765
R12735 VSS.n2113 VSS.n2112 0.2765
R12736 VSS.n2151 VSS.n2150 0.2765
R12737 VSS.n443 VSS.n442 0.26975
R12738 VSS.n686 VSS.n685 0.269
R12739 VSS.n2138 VSS.n2137 0.269
R12740 VSS.n839 VSS.n838 0.26825
R12741 VSS.n1990 VSS.n1989 0.26525
R12742 VSS.n2348 VSS.n89 0.2645
R12743 VSS.n1905 VSS.n1904 0.2645
R12744 VSS.n2174 VSS.n2173 0.2645
R12745 VSS.n500 VSS.n405 0.2645
R12746 VSS.n120 VSS.n119 0.263882
R12747 VSS.n149 VSS.n148 0.263882
R12748 VSS.n178 VSS.n177 0.263882
R12749 VSS.n207 VSS.n206 0.263882
R12750 VSS.n236 VSS.n235 0.263882
R12751 VSS.n291 VSS.n290 0.263882
R12752 VSS.n327 VSS.n326 0.263882
R12753 VSS.n958 VSS.n957 0.26375
R12754 VSS.n943 VSS.n942 0.26375
R12755 VSS.n678 VSS.n677 0.26375
R12756 VSS.n960 VSS.n959 0.263
R12757 VSS.n2407 VSS.n2406 0.2615
R12758 VSS.n736 VSS.n735 0.26
R12759 VSS.n2143 VSS.n2142 0.25775
R12760 VSS.n2249 VSS.n2248 0.2555
R12761 VSS.n964 VSS.n963 0.2555
R12762 VSS.n2216 VSS.n2215 0.2555
R12763 VSS.n1906 VSS.n1905 0.25475
R12764 VSS.n2058 VSS.n2057 0.25475
R12765 VSS.n698 VSS.n697 0.25475
R12766 VSS.n454 VSS.n425 0.25475
R12767 VSS.n1916 VSS.n1915 0.25325
R12768 VSS.n2256 VSS.n2255 0.2525
R12769 VSS.n2258 VSS.n2257 0.2525
R12770 VSS.n2260 VSS.n2259 0.2525
R12771 VSS.n2262 VSS.n2261 0.2525
R12772 VSS.n2264 VSS.n2263 0.2525
R12773 VSS.n2266 VSS.n2265 0.2525
R12774 VSS.n2280 VSS.n2279 0.2525
R12775 VSS.n2278 VSS.n2277 0.2525
R12776 VSS.n2276 VSS.n2275 0.2525
R12777 VSS.n2274 VSS.n2273 0.2525
R12778 VSS.n2272 VSS.n2271 0.2525
R12779 VSS.n2270 VSS.n2269 0.2525
R12780 VSS.n2268 VSS.n93 0.2525
R12781 VSS.n2311 VSS.n2310 0.2525
R12782 VSS.n2307 VSS.n2306 0.2525
R12783 VSS.n2305 VSS.n2304 0.2525
R12784 VSS.n2303 VSS.n2302 0.2525
R12785 VSS.n2301 VSS.n2300 0.2525
R12786 VSS.n2299 VSS.n2298 0.2525
R12787 VSS.n2297 VSS.n2296 0.2525
R12788 VSS.n2295 VSS.n2294 0.2525
R12789 VSS.n2293 VSS.n2292 0.2525
R12790 VSS.n2289 VSS.n2288 0.2525
R12791 VSS.n2287 VSS.n2286 0.2525
R12792 VSS.n2285 VSS.n2284 0.2525
R12793 VSS.n2283 VSS.n2282 0.2525
R12794 VSS.n2353 VSS.n2352 0.2525
R12795 VSS.n2355 VSS.n2354 0.2525
R12796 VSS.n2357 VSS.n2356 0.2525
R12797 VSS.n2361 VSS.n2360 0.2525
R12798 VSS.n2363 VSS.n2362 0.2525
R12799 VSS.n2365 VSS.n2364 0.2525
R12800 VSS.n2367 VSS.n2366 0.2525
R12801 VSS.n2369 VSS.n2368 0.2525
R12802 VSS.n2371 VSS.n2370 0.2525
R12803 VSS.n2373 VSS.n2372 0.2525
R12804 VSS.n2375 VSS.n2374 0.2525
R12805 VSS.n2380 VSS.n2379 0.2525
R12806 VSS.n2378 VSS.n2377 0.2525
R12807 VSS.n2402 VSS.n2401 0.2525
R12808 VSS.n2400 VSS.n2399 0.2525
R12809 VSS.n2398 VSS.n2397 0.2525
R12810 VSS.n2396 VSS.n2395 0.2525
R12811 VSS.n2394 VSS.n2393 0.2525
R12812 VSS.n1142 VSS.n1141 0.2525
R12813 VSS.n1140 VSS.n1139 0.2525
R12814 VSS.n1138 VSS.n1137 0.2525
R12815 VSS.n1136 VSS.n1135 0.2525
R12816 VSS.n1134 VSS.n1133 0.2525
R12817 VSS.n1132 VSS.n1131 0.2525
R12818 VSS.n1128 VSS.n1127 0.2525
R12819 VSS.n1126 VSS.n1125 0.2525
R12820 VSS.n1124 VSS.n1123 0.2525
R12821 VSS.n1122 VSS.n1121 0.2525
R12822 VSS.n1120 VSS.n1119 0.2525
R12823 VSS.n1118 VSS.n1117 0.2525
R12824 VSS.n1116 VSS.n1115 0.2525
R12825 VSS.n1113 VSS.n1112 0.2525
R12826 VSS.n1109 VSS.n1108 0.2525
R12827 VSS.n1107 VSS.n1106 0.2525
R12828 VSS.n1105 VSS.n1104 0.2525
R12829 VSS.n1103 VSS.n1102 0.2525
R12830 VSS.n1101 VSS.n1100 0.2525
R12831 VSS.n1099 VSS.n1098 0.2525
R12832 VSS.n1097 VSS.n1096 0.2525
R12833 VSS.n1095 VSS.n1094 0.2525
R12834 VSS.n1091 VSS.n1090 0.2525
R12835 VSS.n1089 VSS.n1088 0.2525
R12836 VSS.n1087 VSS.n1086 0.2525
R12837 VSS.n1085 VSS.n1084 0.2525
R12838 VSS.n1080 VSS.n1079 0.2525
R12839 VSS.n1078 VSS.n1077 0.2525
R12840 VSS.n1076 VSS.n1075 0.2525
R12841 VSS.n1070 VSS.n1069 0.2525
R12842 VSS.n1068 VSS.n1067 0.2525
R12843 VSS.n1066 VSS.n1065 0.2525
R12844 VSS.n1064 VSS.n1063 0.2525
R12845 VSS.n1062 VSS.n1061 0.2525
R12846 VSS.n1060 VSS.n1059 0.2525
R12847 VSS.n1058 VSS.n1057 0.2525
R12848 VSS.n1628 VSS.n1627 0.2525
R12849 VSS.n1630 VSS.n1629 0.2525
R12850 VSS.n1632 VSS.n1631 0.2525
R12851 VSS.n1634 VSS.n1633 0.2525
R12852 VSS.n1636 VSS.n1635 0.2525
R12853 VSS.n1638 VSS.n1637 0.2525
R12854 VSS.n1642 VSS.n1641 0.2525
R12855 VSS.n1644 VSS.n1643 0.2525
R12856 VSS.n1646 VSS.n1645 0.2525
R12857 VSS.n1648 VSS.n1647 0.2525
R12858 VSS.n1650 VSS.n1649 0.2525
R12859 VSS.n1652 VSS.n1651 0.2525
R12860 VSS.n1654 VSS.n1653 0.2525
R12861 VSS.n1658 VSS.n1657 0.2525
R12862 VSS.n1662 VSS.n1661 0.2525
R12863 VSS.n1664 VSS.n1663 0.2525
R12864 VSS.n1666 VSS.n1665 0.2525
R12865 VSS.n1668 VSS.n1667 0.2525
R12866 VSS.n1670 VSS.n1669 0.2525
R12867 VSS.n1672 VSS.n1671 0.2525
R12868 VSS.n1674 VSS.n1673 0.2525
R12869 VSS.n1676 VSS.n1675 0.2525
R12870 VSS.n1680 VSS.n1679 0.2525
R12871 VSS.n1682 VSS.n1681 0.2525
R12872 VSS.n1684 VSS.n1683 0.2525
R12873 VSS.n1686 VSS.n1685 0.2525
R12874 VSS.n1691 VSS.n1690 0.2525
R12875 VSS.n1693 VSS.n1692 0.2525
R12876 VSS.n1695 VSS.n1694 0.2525
R12877 VSS.n1710 VSS.n1709 0.2525
R12878 VSS.n1618 VSS.n1617 0.2525
R12879 VSS.n1616 VSS.n1615 0.2525
R12880 VSS.n1614 VSS.n1613 0.2525
R12881 VSS.n1612 VSS.n1611 0.2525
R12882 VSS.n1610 VSS.n1609 0.2525
R12883 VSS.n1608 VSS.n1607 0.2525
R12884 VSS.n1604 VSS.n1603 0.2525
R12885 VSS.n1602 VSS.n1601 0.2525
R12886 VSS.n1600 VSS.n1599 0.2525
R12887 VSS.n1598 VSS.n1597 0.2525
R12888 VSS.n1596 VSS.n1595 0.2525
R12889 VSS.n1594 VSS.n1593 0.2525
R12890 VSS.n1592 VSS.n1591 0.2525
R12891 VSS.n1589 VSS.n1588 0.2525
R12892 VSS.n1585 VSS.n1584 0.2525
R12893 VSS.n1583 VSS.n1582 0.2525
R12894 VSS.n1581 VSS.n1580 0.2525
R12895 VSS.n1579 VSS.n1578 0.2525
R12896 VSS.n1577 VSS.n1576 0.2525
R12897 VSS.n1575 VSS.n1574 0.2525
R12898 VSS.n1573 VSS.n1572 0.2525
R12899 VSS.n1571 VSS.n1570 0.2525
R12900 VSS.n1175 VSS.n1174 0.2525
R12901 VSS.n1173 VSS.n1172 0.2525
R12902 VSS.n1171 VSS.n1170 0.2525
R12903 VSS.n1169 VSS.n1168 0.2525
R12904 VSS.n1167 VSS.n1166 0.2525
R12905 VSS.n1165 VSS.n1164 0.2525
R12906 VSS.n1161 VSS.n1160 0.2525
R12907 VSS.n1159 VSS.n1158 0.2525
R12908 VSS.n1157 VSS.n1156 0.2525
R12909 VSS.n1155 VSS.n1154 0.2525
R12910 VSS.n1153 VSS.n1152 0.2525
R12911 VSS.n1151 VSS.n1150 0.2525
R12912 VSS.n1149 VSS.n911 0.2525
R12913 VSS.n1798 VSS.n1797 0.2525
R12914 VSS.n1792 VSS.n1791 0.2525
R12915 VSS.n1790 VSS.n1789 0.2525
R12916 VSS.n1788 VSS.n1787 0.2525
R12917 VSS.n1786 VSS.n1785 0.2525
R12918 VSS.n1784 VSS.n1783 0.2525
R12919 VSS.n1782 VSS.n1781 0.2525
R12920 VSS.n1780 VSS.n1779 0.2525
R12921 VSS.n1205 VSS.n1204 0.2525
R12922 VSS.n1203 VSS.n1202 0.2525
R12923 VSS.n1201 VSS.n1200 0.2525
R12924 VSS.n1199 VSS.n1198 0.2525
R12925 VSS.n1197 VSS.n1196 0.2525
R12926 VSS.n1195 VSS.n1194 0.2525
R12927 VSS.n1191 VSS.n1190 0.2525
R12928 VSS.n1189 VSS.n1188 0.2525
R12929 VSS.n1187 VSS.n1186 0.2525
R12930 VSS.n1185 VSS.n1184 0.2525
R12931 VSS.n1183 VSS.n1182 0.2525
R12932 VSS.n1181 VSS.n1180 0.2525
R12933 VSS.n1179 VSS.n909 0.2525
R12934 VSS.n1804 VSS.n1803 0.2525
R12935 VSS.n1808 VSS.n1807 0.2525
R12936 VSS.n1810 VSS.n1809 0.2525
R12937 VSS.n1812 VSS.n1811 0.2525
R12938 VSS.n1814 VSS.n1813 0.2525
R12939 VSS.n1816 VSS.n1815 0.2525
R12940 VSS.n1818 VSS.n1817 0.2525
R12941 VSS.n1820 VSS.n1819 0.2525
R12942 VSS.n1822 VSS.n1821 0.2525
R12943 VSS.n1826 VSS.n1825 0.2525
R12944 VSS.n1828 VSS.n1827 0.2525
R12945 VSS.n1870 VSS.n1869 0.2525
R12946 VSS.n1265 VSS.n1264 0.2525
R12947 VSS.n1263 VSS.n1262 0.2525
R12948 VSS.n1261 VSS.n1260 0.2525
R12949 VSS.n1259 VSS.n1258 0.2525
R12950 VSS.n1257 VSS.n1256 0.2525
R12951 VSS.n1255 VSS.n1254 0.2525
R12952 VSS.n1251 VSS.n1250 0.2525
R12953 VSS.n1249 VSS.n1248 0.2525
R12954 VSS.n1247 VSS.n1246 0.2525
R12955 VSS.n1245 VSS.n1244 0.2525
R12956 VSS.n1243 VSS.n1242 0.2525
R12957 VSS.n1241 VSS.n1240 0.2525
R12958 VSS.n1239 VSS.n1238 0.2525
R12959 VSS.n1236 VSS.n1235 0.2525
R12960 VSS.n1232 VSS.n1231 0.2525
R12961 VSS.n1230 VSS.n1229 0.2525
R12962 VSS.n1228 VSS.n1227 0.2525
R12963 VSS.n1226 VSS.n1225 0.2525
R12964 VSS.n1224 VSS.n1223 0.2525
R12965 VSS.n1222 VSS.n1221 0.2525
R12966 VSS.n1220 VSS.n1219 0.2525
R12967 VSS.n1218 VSS.n1217 0.2525
R12968 VSS.n1295 VSS.n1294 0.2525
R12969 VSS.n1293 VSS.n1292 0.2525
R12970 VSS.n1291 VSS.n1290 0.2525
R12971 VSS.n1289 VSS.n1288 0.2525
R12972 VSS.n1287 VSS.n1286 0.2525
R12973 VSS.n1285 VSS.n1284 0.2525
R12974 VSS.n1281 VSS.n1280 0.2525
R12975 VSS.n1279 VSS.n1278 0.2525
R12976 VSS.n1277 VSS.n1276 0.2525
R12977 VSS.n1275 VSS.n1274 0.2525
R12978 VSS.n1273 VSS.n1272 0.2525
R12979 VSS.n1271 VSS.n1270 0.2525
R12980 VSS.n1269 VSS.n780 0.2525
R12981 VSS.n1941 VSS.n1940 0.2525
R12982 VSS.n1935 VSS.n1934 0.2525
R12983 VSS.n1933 VSS.n1932 0.2525
R12984 VSS.n1931 VSS.n1930 0.2525
R12985 VSS.n1929 VSS.n1928 0.2525
R12986 VSS.n1927 VSS.n1926 0.2525
R12987 VSS.n1925 VSS.n1924 0.2525
R12988 VSS.n1923 VSS.n1922 0.2525
R12989 VSS.n1325 VSS.n1324 0.2525
R12990 VSS.n1323 VSS.n1322 0.2525
R12991 VSS.n1321 VSS.n1320 0.2525
R12992 VSS.n1319 VSS.n1318 0.2525
R12993 VSS.n1317 VSS.n1316 0.2525
R12994 VSS.n1315 VSS.n1314 0.2525
R12995 VSS.n1311 VSS.n1310 0.2525
R12996 VSS.n1309 VSS.n1308 0.2525
R12997 VSS.n1307 VSS.n1306 0.2525
R12998 VSS.n1305 VSS.n1304 0.2525
R12999 VSS.n1303 VSS.n1302 0.2525
R13000 VSS.n1301 VSS.n1300 0.2525
R13001 VSS.n1299 VSS.n778 0.2525
R13002 VSS.n1947 VSS.n1946 0.2525
R13003 VSS.n1953 VSS.n1952 0.2525
R13004 VSS.n1955 VSS.n1954 0.2525
R13005 VSS.n1957 VSS.n1956 0.2525
R13006 VSS.n1975 VSS.n1974 0.2525
R13007 VSS.n1992 VSS.n1991 0.2525
R13008 VSS.n1396 VSS.n1395 0.2525
R13009 VSS.n1394 VSS.n1393 0.2525
R13010 VSS.n1392 VSS.n1391 0.2525
R13011 VSS.n1390 VSS.n1389 0.2525
R13012 VSS.n1388 VSS.n1387 0.2525
R13013 VSS.n1386 VSS.n1385 0.2525
R13014 VSS.n1362 VSS.n1361 0.2525
R13015 VSS.n1344 VSS.n1343 0.2525
R13016 VSS.n1426 VSS.n1425 0.2525
R13017 VSS.n1424 VSS.n1423 0.2525
R13018 VSS.n1422 VSS.n1421 0.2525
R13019 VSS.n1420 VSS.n1419 0.2525
R13020 VSS.n1418 VSS.n1417 0.2525
R13021 VSS.n1416 VSS.n1415 0.2525
R13022 VSS.n1412 VSS.n1411 0.2525
R13023 VSS.n1410 VSS.n1409 0.2525
R13024 VSS.n1408 VSS.n1407 0.2525
R13025 VSS.n1406 VSS.n1405 0.2525
R13026 VSS.n1404 VSS.n1403 0.2525
R13027 VSS.n1402 VSS.n1401 0.2525
R13028 VSS.n1400 VSS.n635 0.2525
R13029 VSS.n2076 VSS.n2075 0.2525
R13030 VSS.n2070 VSS.n2069 0.2525
R13031 VSS.n2068 VSS.n2067 0.2525
R13032 VSS.n2066 VSS.n2065 0.2525
R13033 VSS.n681 VSS.n680 0.2525
R13034 VSS.n679 VSS.n678 0.2525
R13035 VSS.n1505 VSS.n1504 0.2525
R13036 VSS.n1503 VSS.n1502 0.2525
R13037 VSS.n1501 VSS.n1500 0.2525
R13038 VSS.n1499 VSS.n1498 0.2525
R13039 VSS.n1497 VSS.n1496 0.2525
R13040 VSS.n1495 VSS.n1494 0.2525
R13041 VSS.n1532 VSS.n1531 0.2525
R13042 VSS.n1530 VSS.n1529 0.2525
R13043 VSS.n448 VSS.n447 0.2525
R13044 VSS.n2082 VSS.n2081 0.2525
R13045 VSS.n2064 VSS.n2063 0.25175
R13046 VSS.n1872 VSS.n1871 0.25025
R13047 VSS.n2057 VSS.n2056 0.25025
R13048 VSS.n1715 VSS.n1714 0.2495
R13049 VSS.n2028 VSS.n2027 0.2465
R13050 VSS.n2017 VSS.n2016 0.24425
R13051 VSS.n1053 VSS.n1052 0.2435
R13052 VSS.n956 VSS.n955 0.2435
R13053 VSS.n1879 VSS.n1878 0.2435
R13054 VSS.n2049 VSS.n2048 0.2435
R13055 VSS.n1878 VSS.n1877 0.24275
R13056 VSS.n1907 VSS.n1906 0.24125
R13057 VSS.n2059 VSS.n2058 0.24125
R13058 VSS.n697 VSS.n696 0.24125
R13059 VSS.n455 VSS.n454 0.24125
R13060 VSS.n2124 VSS.n2123 0.24125
R13061 VSS.n1832 VSS.n1831 0.2405
R13062 VSS.n1535 VSS.n1534 0.23975
R13063 VSS.n2137 VSS.n2136 0.239
R13064 VSS.n1753 VSS.n1752 0.23825
R13065 VSS.n600 VSS.n599 0.2375
R13066 VSS.n2169 VSS.n2168 0.23675
R13067 VSS.n941 VSS.n940 0.23375
R13068 VSS.n885 VSS.n884 0.23375
R13069 VSS.n823 VSS.n822 0.23375
R13070 VSS.n1360 VSS.n1359 0.23375
R13071 VSS.n739 VSS.n738 0.23375
R13072 VSS.n677 VSS.n676 0.23375
R13073 VSS.n1486 VSS.n1485 0.23375
R13074 VSS.n2168 VSS.n2167 0.23375
R13075 VSS.n562 VSS.n561 0.23375
R13076 VSS.n1527 VSS.n1526 0.23375
R13077 VSS.n1989 VSS.n1988 0.23075
R13078 VSS.n1001 VSS.n1000 0.2285
R13079 VSS.n1836 VSS.n1835 0.2285
R13080 VSS.n812 VSS.n811 0.2285
R13081 VSS.n2039 VSS.n2038 0.2285
R13082 VSS.n666 VSS.n665 0.2285
R13083 VSS.n573 VSS.n572 0.2285
R13084 VSS.n1436 VSS.n1435 0.2285
R13085 VSS.n1434 VSS.n1433 0.2285
R13086 VSS.n1700 VSS.n1699 0.2255
R13087 VSS.n1702 VSS.n1701 0.2255
R13088 VSS.n1704 VSS.n1703 0.2255
R13089 VSS.n1706 VSS.n1705 0.2255
R13090 VSS.n1708 VSS.n1707 0.2255
R13091 VSS.n848 VSS.n847 0.2255
R13092 VSS.n1982 VSS.n1981 0.2255
R13093 VSS.n1342 VSS.n1341 0.2255
R13094 VSS.n2061 VSS.n2060 0.22325
R13095 VSS.n2158 VSS.n2157 0.22325
R13096 VSS.n2182 VSS.n2181 0.22325
R13097 VSS.n1047 VSS.n1046 0.2225
R13098 VSS.n1715 VSS.n1711 0.2225
R13099 VSS.n1850 VSS.n1849 0.2225
R13100 VSS.n824 VSS.n823 0.2225
R13101 VSS.n1993 VSS.n1992 0.2225
R13102 VSS.n2042 VSS.n2041 0.2225
R13103 VSS.n1472 VSS.n1471 0.2225
R13104 VSS.n457 VSS.n452 0.2225
R13105 VSS.n121 VSS.n110 0.220767
R13106 VSS.n150 VSS.n139 0.220767
R13107 VSS.n179 VSS.n168 0.220767
R13108 VSS.n208 VSS.n197 0.220767
R13109 VSS.n237 VSS.n226 0.220767
R13110 VSS.n299 VSS.n255 0.220767
R13111 VSS.n328 VSS.n317 0.220767
R13112 VSS.n2464 VSS.n2463 0.220767
R13113 VSS.n2198 VSS.n2197 0.2195
R13114 VSS.n742 VSS.n741 0.218
R13115 VSS.n586 VSS.n585 0.2165
R13116 VSS.n1883 VSS.n1882 0.21425
R13117 VSS.n1912 VSS.n1911 0.2135
R13118 VSS.n1972 VSS.n1971 0.2135
R13119 VSS.n558 VSS.n557 0.2075
R13120 VSS.n439 VSS.n404 0.2075
R13121 VSS.n836 VSS.n835 0.2045
R13122 VSS.n2014 VSS.n2013 0.20375
R13123 VSS.n2100 VSS.n2099 0.20375
R13124 VSS.n2141 VSS.n2140 0.20225
R13125 VSS.n2314 VSS.n91 0.2015
R13126 VSS.n1847 VSS.n1846 0.2015
R13127 VSS.n833 VSS.n832 0.2015
R13128 VSS.n684 VSS.n683 0.2015
R13129 VSS.n1541 VSS.n1540 0.2015
R13130 VSS.n966 VSS.n965 0.20075
R13131 VSS.n1759 VSS.n1758 0.1985
R13132 VSS.n743 VSS.n742 0.1985
R13133 VSS.n1441 VSS.n1440 0.1985
R13134 VSS.n2196 VSS.n2195 0.19775
R13135 VSS.n1892 VSS.n1891 0.1955
R13136 VSS.n1353 VSS.n1352 0.1955
R13137 VSS.n1351 VSS.n1350 0.1955
R13138 VSS.n2054 VSS.n2053 0.1955
R13139 VSS.n703 VSS.n702 0.1955
R13140 VSS.n2114 VSS.n2113 0.1955
R13141 VSS.n700 VSS.n699 0.194
R13142 VSS.n1959 VSS.n1958 0.1925
R13143 VSS.n1961 VSS.n1960 0.1925
R13144 VSS.n1963 VSS.n1962 0.1925
R13145 VSS.n2152 VSS.n603 0.191
R13146 VSS.n589 VSS.n588 0.19025
R13147 VSS.n696 VSS.n695 0.18875
R13148 VSS.n962 VSS.n961 0.18725
R13149 VSS.n1537 VSS.n1536 0.18725
R13150 VSS.n594 VSS.n593 0.18725
R13151 VSS.n2542 VSS.n2541 0.185
R13152 VSS.n1897 VSS.n1896 0.18425
R13153 VSS.n596 VSS.n595 0.18425
R13154 VSS.n2019 VSS.n2018 0.18275
R13155 VSS.n2118 VSS.n2117 0.18125
R13156 VSS.n2350 VSS.n87 0.1805
R13157 VSS.n1083 VSS.n1082 0.1805
R13158 VSS.n1688 VSS.n1687 0.1805
R13159 VSS.n1764 VSS.n971 0.1805
R13160 VSS VSS.n0 0.1788
R13161 VSS.n2170 VSS.n2169 0.17825
R13162 VSS.n2404 VSS.n2403 0.1775
R13163 VSS.n441 VSS.n440 0.176
R13164 VSS.n2528 VSS.n2525 0.17375
R13165 VSS.n2171 VSS.n2170 0.173
R13166 VSS.n2167 VSS.n2166 0.1715
R13167 VSS.n1873 VSS.n1872 0.17075
R13168 VSS.n559 VSS.n558 0.17075
R13169 VSS.n2188 VSS.n2187 0.17075
R13170 VSS.n1903 VSS.n1902 0.17
R13171 VSS.n1044 VSS.n1043 0.1685
R13172 VSS.n1005 VSS.n1004 0.1685
R13173 VSS.n999 VSS.n998 0.1685
R13174 VSS.n998 VSS.n997 0.1685
R13175 VSS.n1776 VSS.n1775 0.1685
R13176 VSS.n1775 VSS.n1774 0.1685
R13177 VSS.n1774 VSS.n1773 0.1685
R13178 VSS.n1773 VSS.n1772 0.1685
R13179 VSS.n1772 VSS.n1771 0.1685
R13180 VSS.n1771 VSS.n1770 0.1685
R13181 VSS.n1770 VSS.n1769 0.1685
R13182 VSS.n1769 VSS.n1768 0.1685
R13183 VSS.n969 VSS.n968 0.1685
R13184 VSS.n817 VSS.n816 0.1685
R13185 VSS.n816 VSS.n815 0.1685
R13186 VSS.n2005 VSS.n2004 0.1685
R13187 VSS.n1381 VSS.n1380 0.1685
R13188 VSS.n1380 VSS.n1379 0.1685
R13189 VSS.n1379 VSS.n1378 0.1685
R13190 VSS.n1378 VSS.n1377 0.1685
R13191 VSS.n1377 VSS.n1376 0.1685
R13192 VSS.n1376 VSS.n1375 0.1685
R13193 VSS.n1375 VSS.n1374 0.1685
R13194 VSS.n1374 VSS.n1373 0.1685
R13195 VSS.n1373 VSS.n1372 0.1685
R13196 VSS.n1372 VSS.n1371 0.1685
R13197 VSS.n1371 VSS.n1370 0.1685
R13198 VSS.n1368 VSS.n1367 0.1685
R13199 VSS.n1367 VSS.n1366 0.1685
R13200 VSS.n671 VSS.n670 0.1685
R13201 VSS.n670 VSS.n669 0.1685
R13202 VSS.n568 VSS.n567 0.1685
R13203 VSS.n569 VSS.n568 0.1685
R13204 VSS.n1540 VSS.n1539 0.1685
R13205 VSS.n1539 VSS.n1538 0.1685
R13206 VSS.n582 VSS.n581 0.1685
R13207 VSS.n581 VSS.n580 0.1685
R13208 VSS.n2214 VSS.n2213 0.1685
R13209 VSS.n891 VSS.n890 0.16625
R13210 VSS.n2189 VSS.n2188 0.16625
R13211 VSS.n834 VSS.n833 0.1655
R13212 VSS.n953 VSS.n952 0.16475
R13213 VSS.n942 VSS.n941 0.16475
R13214 VSS.n832 VSS.n831 0.16475
R13215 VSS.n688 VSS.n687 0.16475
R13216 VSS.n1848 VSS.n1847 0.1625
R13217 VSS.n274 VSS.n272 0.161
R13218 VSS.n2025 VSS.n748 0.161
R13219 VSS.n279 VSS.n277 0.1605
R13220 VSS.n281 VSS.n279 0.1605
R13221 VSS.n270 VSS.n268 0.1605
R13222 VSS.n272 VSS.n270 0.1605
R13223 VSS.n2552 VSS.n2551 0.159626
R13224 VSS.n1483 VSS.n1482 0.1595
R13225 VSS.n952 VSS.n951 0.15875
R13226 VSS.n829 VSS.n828 0.15875
R13227 VSS.n2520 VSS.n2518 0.158515
R13228 VSS.n283 VSS.n281 0.1585
R13229 VSS.n1764 VSS.n1763 0.1565
R13230 VSS.n1767 VSS.n969 0.1565
R13231 VSS.n1898 VSS.n1897 0.15575
R13232 VSS.n2119 VSS.n2118 0.15575
R13233 VSS.n845 VSS.n844 0.15425
R13234 VSS.n2020 VSS.n2019 0.15425
R13235 VSS.n2148 VSS.n2147 0.1535
R13236 VSS.n748 VSS.n747 0.152
R13237 VSS.n1538 VSS.n1537 0.14975
R13238 VSS.n1841 VSS.n1840 0.14825
R13239 VSS.n1890 VSS.n1889 0.14825
R13240 VSS.n695 VSS.n694 0.14825
R13241 VSS.n1470 VSS.n1469 0.14825
R13242 VSS.n590 VSS.n589 0.14675
R13243 VSS.n1876 VSS.n1875 0.146
R13244 VSS.n1960 VSS.n1959 0.1445
R13245 VSS.n1962 VSS.n1961 0.1445
R13246 VSS.n1964 VSS.n1963 0.1445
R13247 VSS.n2045 VSS.n2044 0.1445
R13248 VSS.n2062 VSS.n2061 0.14375
R13249 VSS.n2497 VSS.n2496 0.143273
R13250 VSS.n1888 VSS.n1887 0.14225
R13251 VSS.n1346 VSS.n1345 0.14225
R13252 VSS.n1758 VSS.n1757 0.1415
R13253 VSS.n1354 VSS.n1353 0.1415
R13254 VSS.n1352 VSS.n1351 0.1415
R13255 VSS.n2080 VSS.n633 0.1415
R13256 VSS.n2509 VSS.n2508 0.141125
R13257 VSS.n122 VSS.n121 0.140132
R13258 VSS.n151 VSS.n150 0.140132
R13259 VSS.n180 VSS.n179 0.140132
R13260 VSS.n209 VSS.n208 0.140132
R13261 VSS.n238 VSS.n237 0.140132
R13262 VSS.n300 VSS.n299 0.140132
R13263 VSS.n329 VSS.n328 0.140132
R13264 VSS.n262 VSS.n259 0.139126
R13265 VSS.n2240 VSS.n2239 0.1385
R13266 VSS.n2318 VSS.n2317 0.1385
R13267 VSS.n2329 VSS.n2326 0.1385
R13268 VSS.n2343 VSS.n2342 0.1385
R13269 VSS.n2334 VSS.n2333 0.1385
R13270 VSS.n2412 VSS.n2411 0.1385
R13271 VSS.n2281 VSS.n2267 0.1385
R13272 VSS.n2309 VSS.n2308 0.1385
R13273 VSS.n2291 VSS.n2290 0.1385
R13274 VSS.n2359 VSS.n2358 0.1385
R13275 VSS.n2381 VSS.n2376 0.1385
R13276 VSS.n2392 VSS.n2391 0.1385
R13277 VSS.n1130 VSS.n1129 0.1385
R13278 VSS.n1111 VSS.n1110 0.1385
R13279 VSS.n1093 VSS.n1092 0.1385
R13280 VSS.n1074 VSS.n1073 0.1385
R13281 VSS.n1640 VSS.n1639 0.1385
R13282 VSS.n1660 VSS.n1659 0.1385
R13283 VSS.n1678 VSS.n1677 0.1385
R13284 VSS.n1697 VSS.n1696 0.1385
R13285 VSS.n1606 VSS.n1605 0.1385
R13286 VSS.n1587 VSS.n1586 0.1385
R13287 VSS.n1569 VSS.n1568 0.1385
R13288 VSS.n1760 VSS.n1759 0.1385
R13289 VSS.n1163 VSS.n1162 0.1385
R13290 VSS.n1796 VSS.n1795 0.1385
R13291 VSS.n1193 VSS.n1192 0.1385
R13292 VSS.n1806 VSS.n1805 0.1385
R13293 VSS.n1824 VSS.n1823 0.1385
R13294 VSS.n1253 VSS.n1252 0.1385
R13295 VSS.n1234 VSS.n1233 0.1385
R13296 VSS.n1216 VSS.n1215 0.1385
R13297 VSS.n1283 VSS.n1282 0.1385
R13298 VSS.n1939 VSS.n1938 0.1385
R13299 VSS.n843 VSS.n842 0.1385
R13300 VSS.n1313 VSS.n1312 0.1385
R13301 VSS.n1949 VSS.n1948 0.1385
R13302 VSS.n1965 VSS.n1964 0.1385
R13303 VSS.n1980 VSS.n1979 0.1385
R13304 VSS.n1384 VSS.n1383 0.1385
R13305 VSS.n1366 VSS.n1365 0.1385
R13306 VSS.n1350 VSS.n1349 0.1385
R13307 VSS.n2030 VSS.n2029 0.1385
R13308 VSS.n1414 VSS.n1413 0.1385
R13309 VSS.n2074 VSS.n2073 0.1385
R13310 VSS.n1493 VSS.n1492 0.1385
R13311 VSS.n457 VSS.n456 0.1385
R13312 VSS.n1442 VSS.n1441 0.1385
R13313 VSS.n2207 VSS.n2206 0.1385
R13314 VSS.n503 VSS.n497 0.1385
R13315 VSS.n515 VSS.n514 0.1385
R13316 VSS.n525 VSS.n523 0.1385
R13317 VSS.n533 VSS.n532 0.1385
R13318 VSS.n2315 VSS.n2314 0.1355
R13319 VSS.n2081 VSS.n2080 0.1355
R13320 VSS.n296 VSS.n259 0.13486
R13321 VSS.n2139 VSS.n2138 0.13475
R13322 VSS.n563 VSS.n562 0.13325
R13323 VSS.n1526 VSS.n1525 0.13325
R13324 VSS.n600 VSS.n425 0.13325
R13325 VSS.n2099 VSS.n2098 0.13325
R13326 VSS.n1469 VSS.n1468 0.13175
R13327 VSS.n556 VSS.n422 0.13175
R13328 VSS.n2179 VSS.n2178 0.13175
R13329 VSS.n2498 VSS.n2497 0.131409
R13330 VSS.n2507 VSS.n2506 0.131409
R13331 VSS.n675 VSS.n674 0.12875
R13332 VSS.n2117 VSS.n2116 0.12875
R13333 VSS.n47 VSS.n46 0.12686
R13334 VSS.n2009 VSS.n2008 0.12125
R13335 VSS.n1522 VSS.n1521 0.12125
R13336 VSS.n2092 VSS.n2091 0.12125
R13337 VSS.n2250 VSS.n358 0.1205
R13338 VSS.n2252 VSS.n95 0.1205
R13339 VSS.n1146 VSS.n1145 0.1205
R13340 VSS.n1624 VSS.n1147 0.1205
R13341 VSS.n1621 VSS.n1563 0.1205
R13342 VSS.n1562 VSS.n1178 0.1205
R13343 VSS.n1561 VSS.n1208 0.1205
R13344 VSS.n1560 VSS.n1268 0.1205
R13345 VSS.n1559 VSS.n1298 0.1205
R13346 VSS.n1558 VSS.n1328 0.1205
R13347 VSS.n1557 VSS.n1399 0.1205
R13348 VSS.n1556 VSS.n1429 0.1205
R13349 VSS.n693 VSS.n692 0.1205
R13350 VSS.n1554 VSS.n1508 0.1205
R13351 VSS.n1553 VSS.n1551 0.1205
R13352 VSS.n587 VSS.n586 0.1205
R13353 VSS.n1555 VSS.n1450 0.1205
R13354 VSS.n2098 VSS.n2097 0.1205
R13355 VSS.n1552 VSS.n373 0.1205
R13356 VSS.n1843 VSS.n1842 0.11825
R13357 VSS.n1849 VSS.n1848 0.1175
R13358 VSS.n1370 VSS.n1369 0.1175
R13359 VSS.n1339 VSS.n706 0.1175
R13360 VSS.n732 VSS.n731 0.1175
R13361 VSS.n2194 VSS.n2193 0.1175
R13362 VSS.n2110 VSS.n2109 0.1175
R13363 VSS.n2152 VSS.n2151 0.1175
R13364 VSS.n946 VSS.n945 0.11675
R13365 VSS.n2097 VSS.n2096 0.11675
R13366 VSS.n126 VSS.n125 0.115978
R13367 VSS.n119 VSS.n118 0.115978
R13368 VSS.n155 VSS.n154 0.115978
R13369 VSS.n148 VSS.n147 0.115978
R13370 VSS.n184 VSS.n183 0.115978
R13371 VSS.n177 VSS.n176 0.115978
R13372 VSS.n213 VSS.n212 0.115978
R13373 VSS.n206 VSS.n205 0.115978
R13374 VSS.n242 VSS.n241 0.115978
R13375 VSS.n235 VSS.n234 0.115978
R13376 VSS.n290 VSS.n289 0.115978
R13377 VSS.n304 VSS.n303 0.115978
R13378 VSS.n333 VSS.n332 0.115978
R13379 VSS.n326 VSS.n325 0.115978
R13380 VSS.n21 VSS.n20 0.1157
R13381 VSS.n46 VSS.n45 0.1157
R13382 VSS.n889 VSS.n888 0.11525
R13383 VSS.n2281 VSS.n2280 0.1145
R13384 VSS.n2308 VSS.n2307 0.1145
R13385 VSS.n2290 VSS.n2289 0.1145
R13386 VSS.n2360 VSS.n2359 0.1145
R13387 VSS.n2381 VSS.n2380 0.1145
R13388 VSS.n2391 VSS.n2390 0.1145
R13389 VSS.n1129 VSS.n1128 0.1145
R13390 VSS.n1110 VSS.n1109 0.1145
R13391 VSS.n1092 VSS.n1091 0.1145
R13392 VSS.n1073 VSS.n1072 0.1145
R13393 VSS.n1046 VSS.n1045 0.1145
R13394 VSS.n1641 VSS.n1640 0.1145
R13395 VSS.n1661 VSS.n1660 0.1145
R13396 VSS.n1679 VSS.n1678 0.1145
R13397 VSS.n1698 VSS.n1697 0.1145
R13398 VSS.n1605 VSS.n1604 0.1145
R13399 VSS.n1586 VSS.n1585 0.1145
R13400 VSS.n1568 VSS.n1567 0.1145
R13401 VSS.n1162 VSS.n1161 0.1145
R13402 VSS.n1795 VSS.n1794 0.1145
R13403 VSS.n940 VSS.n939 0.1145
R13404 VSS.n1192 VSS.n1191 0.1145
R13405 VSS.n1807 VSS.n1806 0.1145
R13406 VSS.n1825 VSS.n1824 0.1145
R13407 VSS.n1252 VSS.n1251 0.1145
R13408 VSS.n1233 VSS.n1232 0.1145
R13409 VSS.n1215 VSS.n1214 0.1145
R13410 VSS.n884 VSS.n883 0.1145
R13411 VSS.n1282 VSS.n1281 0.1145
R13412 VSS.n1938 VSS.n1937 0.1145
R13413 VSS.n1312 VSS.n1311 0.1145
R13414 VSS.n1950 VSS.n1949 0.1145
R13415 VSS.n1383 VSS.n1382 0.1145
R13416 VSS.n2043 VSS.n2042 0.1145
R13417 VSS.n1413 VSS.n1412 0.1145
R13418 VSS.n2073 VSS.n2072 0.1145
R13419 VSS.n1701 VSS.n1700 0.1115
R13420 VSS.n1703 VSS.n1702 0.1115
R13421 VSS.n1705 VSS.n1704 0.1115
R13422 VSS.n1707 VSS.n1706 0.1115
R13423 VSS.n1709 VSS.n1708 0.1115
R13424 VSS.n1211 VSS.n1210 0.1115
R13425 VSS.n847 VSS.n846 0.1115
R13426 VSS.n1343 VSS.n1342 0.1115
R13427 VSS.n1341 VSS.n1340 0.1115
R13428 VSS.n1347 VSS.n1346 0.11075
R13429 VSS.n967 VSS.n966 0.10925
R13430 VSS.n1213 VSS.n1212 0.10925
R13431 VSS.n2197 VSS.n2196 0.10925
R13432 VSS.n447 VSS.n446 0.10925
R13433 VSS.n2086 VSS.n2085 0.10925
R13434 VSS.n488 VSS.n487 0.10925
R13435 VSS.n2414 VSS.n2413 0.1085
R13436 VSS.n1043 VSS.n1042 0.1085
R13437 VSS.n1006 VSS.n1005 0.1085
R13438 VSS.n1000 VSS.n999 0.1085
R13439 VSS.n934 VSS.n933 0.1085
R13440 VSS.n1893 VSS.n1892 0.1085
R13441 VSS.n878 VSS.n877 0.1085
R13442 VSS.n1917 VSS.n1916 0.1085
R13443 VSS.n811 VSS.n810 0.1085
R13444 VSS.n1986 VSS.n1985 0.1085
R13445 VSS.n1340 VSS.n1339 0.1085
R13446 VSS.n2038 VSS.n2037 0.1085
R13447 VSS.n665 VSS.n664 0.1085
R13448 VSS.n574 VSS.n573 0.1085
R13449 VSS.n1437 VSS.n1436 0.1085
R13450 VSS.n1435 VSS.n1434 0.1085
R13451 VSS.n125 VSS.n124 0.106382
R13452 VSS.n118 VSS.n117 0.106382
R13453 VSS.n154 VSS.n153 0.106382
R13454 VSS.n147 VSS.n146 0.106382
R13455 VSS.n183 VSS.n182 0.106382
R13456 VSS.n176 VSS.n175 0.106382
R13457 VSS.n212 VSS.n211 0.106382
R13458 VSS.n205 VSS.n204 0.106382
R13459 VSS.n241 VSS.n240 0.106382
R13460 VSS.n234 VSS.n233 0.106382
R13461 VSS.n289 VSS.n288 0.106382
R13462 VSS.n303 VSS.n302 0.106382
R13463 VSS.n332 VSS.n331 0.106382
R13464 VSS.n325 VSS.n324 0.106382
R13465 VSS.n822 VSS.n821 0.10625
R13466 VSS.n123 VSS.n122 0.106051
R13467 VSS.n116 VSS.n115 0.106051
R13468 VSS.n152 VSS.n151 0.106051
R13469 VSS.n145 VSS.n144 0.106051
R13470 VSS.n181 VSS.n180 0.106051
R13471 VSS.n174 VSS.n173 0.106051
R13472 VSS.n210 VSS.n209 0.106051
R13473 VSS.n203 VSS.n202 0.106051
R13474 VSS.n239 VSS.n238 0.106051
R13475 VSS.n232 VSS.n231 0.106051
R13476 VSS.n287 VSS.n286 0.106051
R13477 VSS.n301 VSS.n300 0.106051
R13478 VSS.n330 VSS.n329 0.106051
R13479 VSS.n323 VSS.n322 0.106051
R13480 VSS.n124 VSS.n123 0.105721
R13481 VSS.n117 VSS.n116 0.105721
R13482 VSS.n153 VSS.n152 0.105721
R13483 VSS.n146 VSS.n145 0.105721
R13484 VSS.n182 VSS.n181 0.105721
R13485 VSS.n175 VSS.n174 0.105721
R13486 VSS.n211 VSS.n210 0.105721
R13487 VSS.n204 VSS.n203 0.105721
R13488 VSS.n240 VSS.n239 0.105721
R13489 VSS.n233 VSS.n232 0.105721
R13490 VSS.n288 VSS.n287 0.105721
R13491 VSS.n302 VSS.n301 0.105721
R13492 VSS.n331 VSS.n330 0.105721
R13493 VSS.n324 VSS.n323 0.105721
R13494 VSS.n689 VSS.n688 0.10475
R13495 VSS.n2013 VSS.n2012 0.10325
R13496 VSS.n1359 VSS.n1358 0.10325
R13497 VSS.n1485 VSS.n1484 0.10325
R13498 VSS.n293 VSS.n291 0.102118
R13499 VSS.n1887 VSS.n1886 0.10175
R13500 VSS.n1754 VSS.n1753 0.09875
R13501 VSS.n2104 VSS.n2103 0.09875
R13502 VSS.n1838 VSS.n1837 0.098
R13503 VSS.n1973 VSS.n1972 0.09725
R13504 VSS.n1534 VSS.n1533 0.09725
R13505 VSS.n2116 VSS.n2115 0.09725
R13506 VSS.n1833 VSS.n1832 0.0965
R13507 VSS.n1911 VSS.n850 0.0965
R13508 VSS.n1492 VSS.n1491 0.09575
R13509 VSS.n456 VSS.n455 0.09575
R13510 VSS.n2105 VSS.n2104 0.095
R13511 VSS.n1052 VSS.n1051 0.0935
R13512 VSS.n1741 VSS.n1014 0.0935
R13513 VSS.n2016 VSS.n2015 0.09275
R13514 VSS.n595 VSS.n594 0.09275
R13515 VSS.n2089 VSS.n2088 0.09275
R13516 VSS.n2508 VSS.n2507 0.0925455
R13517 VSS.n954 VSS.n953 0.09125
R13518 VSS.n22 VSS.n21 0.09086
R13519 VSS.n2029 VSS.n2028 0.0905
R13520 VSS.n339 VSS.n126 0.0878529
R13521 VSS.n338 VSS.n155 0.0878529
R13522 VSS.n337 VSS.n184 0.0878529
R13523 VSS.n336 VSS.n213 0.0878529
R13524 VSS.n335 VSS.n242 0.0878529
R13525 VSS.n334 VSS.n333 0.0878529
R13526 VSS.n699 VSS.n698 0.08675
R13527 VSS.n830 VSS.n829 0.08525
R13528 VSS.n685 VSS.n684 0.08525
R13529 VSS.n2255 VSS.n2254 0.0845
R13530 VSS.n2257 VSS.n2256 0.0845
R13531 VSS.n2259 VSS.n2258 0.0845
R13532 VSS.n2261 VSS.n2260 0.0845
R13533 VSS.n2263 VSS.n2262 0.0845
R13534 VSS.n2265 VSS.n2264 0.0845
R13535 VSS.n2267 VSS.n2266 0.0845
R13536 VSS.n2279 VSS.n2278 0.0845
R13537 VSS.n2277 VSS.n2276 0.0845
R13538 VSS.n2275 VSS.n2274 0.0845
R13539 VSS.n2273 VSS.n2272 0.0845
R13540 VSS.n2271 VSS.n2270 0.0845
R13541 VSS.n2269 VSS.n2268 0.0845
R13542 VSS.n2310 VSS.n2309 0.0845
R13543 VSS.n2306 VSS.n2305 0.0845
R13544 VSS.n2304 VSS.n2303 0.0845
R13545 VSS.n2302 VSS.n2301 0.0845
R13546 VSS.n2300 VSS.n2299 0.0845
R13547 VSS.n2298 VSS.n2297 0.0845
R13548 VSS.n2296 VSS.n2295 0.0845
R13549 VSS.n2294 VSS.n2293 0.0845
R13550 VSS.n2292 VSS.n2291 0.0845
R13551 VSS.n2288 VSS.n2287 0.0845
R13552 VSS.n2286 VSS.n2285 0.0845
R13553 VSS.n2284 VSS.n2283 0.0845
R13554 VSS.n2282 VSS.n87 0.0845
R13555 VSS.n2352 VSS.n2351 0.0845
R13556 VSS.n2354 VSS.n2353 0.0845
R13557 VSS.n2356 VSS.n2355 0.0845
R13558 VSS.n2358 VSS.n2357 0.0845
R13559 VSS.n2362 VSS.n2361 0.0845
R13560 VSS.n2364 VSS.n2363 0.0845
R13561 VSS.n2366 VSS.n2365 0.0845
R13562 VSS.n2368 VSS.n2367 0.0845
R13563 VSS.n2370 VSS.n2369 0.0845
R13564 VSS.n2372 VSS.n2371 0.0845
R13565 VSS.n2374 VSS.n2373 0.0845
R13566 VSS.n2376 VSS.n2375 0.0845
R13567 VSS.n2379 VSS.n2378 0.0845
R13568 VSS.n2377 VSS.n86 0.0845
R13569 VSS.n2403 VSS.n2402 0.0845
R13570 VSS.n2401 VSS.n2400 0.0845
R13571 VSS.n2399 VSS.n2398 0.0845
R13572 VSS.n2397 VSS.n2396 0.0845
R13573 VSS.n2395 VSS.n2394 0.0845
R13574 VSS.n2393 VSS.n2392 0.0845
R13575 VSS.n1143 VSS.n1142 0.0845
R13576 VSS.n1141 VSS.n1140 0.0845
R13577 VSS.n1139 VSS.n1138 0.0845
R13578 VSS.n1137 VSS.n1136 0.0845
R13579 VSS.n1135 VSS.n1134 0.0845
R13580 VSS.n1133 VSS.n1132 0.0845
R13581 VSS.n1131 VSS.n1130 0.0845
R13582 VSS.n1127 VSS.n1126 0.0845
R13583 VSS.n1125 VSS.n1124 0.0845
R13584 VSS.n1123 VSS.n1122 0.0845
R13585 VSS.n1121 VSS.n1120 0.0845
R13586 VSS.n1119 VSS.n1118 0.0845
R13587 VSS.n1117 VSS.n1116 0.0845
R13588 VSS.n1112 VSS.n1111 0.0845
R13589 VSS.n1108 VSS.n1107 0.0845
R13590 VSS.n1106 VSS.n1105 0.0845
R13591 VSS.n1104 VSS.n1103 0.0845
R13592 VSS.n1102 VSS.n1101 0.0845
R13593 VSS.n1100 VSS.n1099 0.0845
R13594 VSS.n1098 VSS.n1097 0.0845
R13595 VSS.n1096 VSS.n1095 0.0845
R13596 VSS.n1094 VSS.n1093 0.0845
R13597 VSS.n1090 VSS.n1089 0.0845
R13598 VSS.n1088 VSS.n1087 0.0845
R13599 VSS.n1086 VSS.n1085 0.0845
R13600 VSS.n1084 VSS.n1083 0.0845
R13601 VSS.n1081 VSS.n1080 0.0845
R13602 VSS.n1079 VSS.n1078 0.0845
R13603 VSS.n1077 VSS.n1076 0.0845
R13604 VSS.n1075 VSS.n1074 0.0845
R13605 VSS.n1071 VSS.n1070 0.0845
R13606 VSS.n1069 VSS.n1068 0.0845
R13607 VSS.n1067 VSS.n1066 0.0845
R13608 VSS.n1065 VSS.n1064 0.0845
R13609 VSS.n1063 VSS.n1062 0.0845
R13610 VSS.n1061 VSS.n1060 0.0845
R13611 VSS.n1059 VSS.n1058 0.0845
R13612 VSS.n1057 VSS.n1056 0.0845
R13613 VSS.n1627 VSS.n1626 0.0845
R13614 VSS.n1629 VSS.n1628 0.0845
R13615 VSS.n1631 VSS.n1630 0.0845
R13616 VSS.n1633 VSS.n1632 0.0845
R13617 VSS.n1635 VSS.n1634 0.0845
R13618 VSS.n1637 VSS.n1636 0.0845
R13619 VSS.n1639 VSS.n1638 0.0845
R13620 VSS.n1643 VSS.n1642 0.0845
R13621 VSS.n1645 VSS.n1644 0.0845
R13622 VSS.n1647 VSS.n1646 0.0845
R13623 VSS.n1649 VSS.n1648 0.0845
R13624 VSS.n1651 VSS.n1650 0.0845
R13625 VSS.n1653 VSS.n1652 0.0845
R13626 VSS.n1659 VSS.n1658 0.0845
R13627 VSS.n1663 VSS.n1662 0.0845
R13628 VSS.n1665 VSS.n1664 0.0845
R13629 VSS.n1667 VSS.n1666 0.0845
R13630 VSS.n1669 VSS.n1668 0.0845
R13631 VSS.n1671 VSS.n1670 0.0845
R13632 VSS.n1673 VSS.n1672 0.0845
R13633 VSS.n1675 VSS.n1674 0.0845
R13634 VSS.n1677 VSS.n1676 0.0845
R13635 VSS.n1681 VSS.n1680 0.0845
R13636 VSS.n1683 VSS.n1682 0.0845
R13637 VSS.n1685 VSS.n1684 0.0845
R13638 VSS.n1687 VSS.n1686 0.0845
R13639 VSS.n1690 VSS.n1689 0.0845
R13640 VSS.n1692 VSS.n1691 0.0845
R13641 VSS.n1694 VSS.n1693 0.0845
R13642 VSS.n1696 VSS.n1695 0.0845
R13643 VSS.n1619 VSS.n1618 0.0845
R13644 VSS.n1617 VSS.n1616 0.0845
R13645 VSS.n1615 VSS.n1614 0.0845
R13646 VSS.n1613 VSS.n1612 0.0845
R13647 VSS.n1611 VSS.n1610 0.0845
R13648 VSS.n1609 VSS.n1608 0.0845
R13649 VSS.n1607 VSS.n1606 0.0845
R13650 VSS.n1603 VSS.n1602 0.0845
R13651 VSS.n1601 VSS.n1600 0.0845
R13652 VSS.n1599 VSS.n1598 0.0845
R13653 VSS.n1597 VSS.n1596 0.0845
R13654 VSS.n1595 VSS.n1594 0.0845
R13655 VSS.n1593 VSS.n1592 0.0845
R13656 VSS.n1588 VSS.n1587 0.0845
R13657 VSS.n1584 VSS.n1583 0.0845
R13658 VSS.n1582 VSS.n1581 0.0845
R13659 VSS.n1580 VSS.n1579 0.0845
R13660 VSS.n1578 VSS.n1577 0.0845
R13661 VSS.n1576 VSS.n1575 0.0845
R13662 VSS.n1574 VSS.n1573 0.0845
R13663 VSS.n1572 VSS.n1571 0.0845
R13664 VSS.n1570 VSS.n1569 0.0845
R13665 VSS.n1176 VSS.n1175 0.0845
R13666 VSS.n1174 VSS.n1173 0.0845
R13667 VSS.n1172 VSS.n1171 0.0845
R13668 VSS.n1170 VSS.n1169 0.0845
R13669 VSS.n1168 VSS.n1167 0.0845
R13670 VSS.n1166 VSS.n1165 0.0845
R13671 VSS.n1164 VSS.n1163 0.0845
R13672 VSS.n1160 VSS.n1159 0.0845
R13673 VSS.n1158 VSS.n1157 0.0845
R13674 VSS.n1156 VSS.n1155 0.0845
R13675 VSS.n1154 VSS.n1153 0.0845
R13676 VSS.n1152 VSS.n1151 0.0845
R13677 VSS.n1150 VSS.n1149 0.0845
R13678 VSS.n1797 VSS.n1796 0.0845
R13679 VSS.n1793 VSS.n1792 0.0845
R13680 VSS.n1791 VSS.n1790 0.0845
R13681 VSS.n1789 VSS.n1788 0.0845
R13682 VSS.n1787 VSS.n1786 0.0845
R13683 VSS.n1785 VSS.n1784 0.0845
R13684 VSS.n1783 VSS.n1782 0.0845
R13685 VSS.n1781 VSS.n1780 0.0845
R13686 VSS.n1779 VSS.n1778 0.0845
R13687 VSS.n1206 VSS.n1205 0.0845
R13688 VSS.n1204 VSS.n1203 0.0845
R13689 VSS.n1202 VSS.n1201 0.0845
R13690 VSS.n1200 VSS.n1199 0.0845
R13691 VSS.n1198 VSS.n1197 0.0845
R13692 VSS.n1196 VSS.n1195 0.0845
R13693 VSS.n1194 VSS.n1193 0.0845
R13694 VSS.n1190 VSS.n1189 0.0845
R13695 VSS.n1188 VSS.n1187 0.0845
R13696 VSS.n1186 VSS.n1185 0.0845
R13697 VSS.n1184 VSS.n1183 0.0845
R13698 VSS.n1182 VSS.n1181 0.0845
R13699 VSS.n1180 VSS.n1179 0.0845
R13700 VSS.n1805 VSS.n1804 0.0845
R13701 VSS.n1809 VSS.n1808 0.0845
R13702 VSS.n1811 VSS.n1810 0.0845
R13703 VSS.n1813 VSS.n1812 0.0845
R13704 VSS.n1815 VSS.n1814 0.0845
R13705 VSS.n1817 VSS.n1816 0.0845
R13706 VSS.n1819 VSS.n1818 0.0845
R13707 VSS.n1821 VSS.n1820 0.0845
R13708 VSS.n1823 VSS.n1822 0.0845
R13709 VSS.n1827 VSS.n1826 0.0845
R13710 VSS.n1882 VSS.n1881 0.0845
R13711 VSS.n1880 VSS.n1879 0.0845
R13712 VSS.n1869 VSS.n1868 0.0845
R13713 VSS.n1266 VSS.n1265 0.0845
R13714 VSS.n1264 VSS.n1263 0.0845
R13715 VSS.n1262 VSS.n1261 0.0845
R13716 VSS.n1260 VSS.n1259 0.0845
R13717 VSS.n1258 VSS.n1257 0.0845
R13718 VSS.n1256 VSS.n1255 0.0845
R13719 VSS.n1254 VSS.n1253 0.0845
R13720 VSS.n1250 VSS.n1249 0.0845
R13721 VSS.n1248 VSS.n1247 0.0845
R13722 VSS.n1246 VSS.n1245 0.0845
R13723 VSS.n1244 VSS.n1243 0.0845
R13724 VSS.n1242 VSS.n1241 0.0845
R13725 VSS.n1240 VSS.n1239 0.0845
R13726 VSS.n1235 VSS.n1234 0.0845
R13727 VSS.n1231 VSS.n1230 0.0845
R13728 VSS.n1229 VSS.n1228 0.0845
R13729 VSS.n1227 VSS.n1226 0.0845
R13730 VSS.n1225 VSS.n1224 0.0845
R13731 VSS.n1223 VSS.n1222 0.0845
R13732 VSS.n1221 VSS.n1220 0.0845
R13733 VSS.n1219 VSS.n1218 0.0845
R13734 VSS.n1217 VSS.n1216 0.0845
R13735 VSS.n1296 VSS.n1295 0.0845
R13736 VSS.n1294 VSS.n1293 0.0845
R13737 VSS.n1292 VSS.n1291 0.0845
R13738 VSS.n1290 VSS.n1289 0.0845
R13739 VSS.n1288 VSS.n1287 0.0845
R13740 VSS.n1286 VSS.n1285 0.0845
R13741 VSS.n1284 VSS.n1283 0.0845
R13742 VSS.n1280 VSS.n1279 0.0845
R13743 VSS.n1278 VSS.n1277 0.0845
R13744 VSS.n1276 VSS.n1275 0.0845
R13745 VSS.n1274 VSS.n1273 0.0845
R13746 VSS.n1272 VSS.n1271 0.0845
R13747 VSS.n1270 VSS.n1269 0.0845
R13748 VSS.n1940 VSS.n1939 0.0845
R13749 VSS.n1936 VSS.n1935 0.0845
R13750 VSS.n1934 VSS.n1933 0.0845
R13751 VSS.n1932 VSS.n1931 0.0845
R13752 VSS.n1930 VSS.n1929 0.0845
R13753 VSS.n1928 VSS.n1927 0.0845
R13754 VSS.n1926 VSS.n1925 0.0845
R13755 VSS.n1924 VSS.n1923 0.0845
R13756 VSS.n1922 VSS.n1921 0.0845
R13757 VSS.n828 VSS.n827 0.0845
R13758 VSS.n826 VSS.n825 0.0845
R13759 VSS.n1326 VSS.n1325 0.0845
R13760 VSS.n1324 VSS.n1323 0.0845
R13761 VSS.n1322 VSS.n1321 0.0845
R13762 VSS.n1320 VSS.n1319 0.0845
R13763 VSS.n1318 VSS.n1317 0.0845
R13764 VSS.n1316 VSS.n1315 0.0845
R13765 VSS.n1314 VSS.n1313 0.0845
R13766 VSS.n1310 VSS.n1309 0.0845
R13767 VSS.n1308 VSS.n1307 0.0845
R13768 VSS.n1306 VSS.n1305 0.0845
R13769 VSS.n1304 VSS.n1303 0.0845
R13770 VSS.n1302 VSS.n1301 0.0845
R13771 VSS.n1300 VSS.n1299 0.0845
R13772 VSS.n1948 VSS.n1947 0.0845
R13773 VSS.n1952 VSS.n1951 0.0845
R13774 VSS.n1954 VSS.n1953 0.0845
R13775 VSS.n1956 VSS.n1955 0.0845
R13776 VSS.n1976 VSS.n1975 0.0845
R13777 VSS.n1991 VSS.n751 0.0845
R13778 VSS.n1397 VSS.n1396 0.0845
R13779 VSS.n1395 VSS.n1394 0.0845
R13780 VSS.n1393 VSS.n1392 0.0845
R13781 VSS.n1391 VSS.n1390 0.0845
R13782 VSS.n1389 VSS.n1388 0.0845
R13783 VSS.n1387 VSS.n1386 0.0845
R13784 VSS.n1385 VSS.n1384 0.0845
R13785 VSS.n1363 VSS.n1362 0.0845
R13786 VSS.n1361 VSS.n1360 0.0845
R13787 VSS.n1345 VSS.n1344 0.0845
R13788 VSS.n1427 VSS.n1426 0.0845
R13789 VSS.n1425 VSS.n1424 0.0845
R13790 VSS.n1423 VSS.n1422 0.0845
R13791 VSS.n1421 VSS.n1420 0.0845
R13792 VSS.n1419 VSS.n1418 0.0845
R13793 VSS.n1417 VSS.n1416 0.0845
R13794 VSS.n1415 VSS.n1414 0.0845
R13795 VSS.n1411 VSS.n1410 0.0845
R13796 VSS.n1409 VSS.n1408 0.0845
R13797 VSS.n1407 VSS.n1406 0.0845
R13798 VSS.n1405 VSS.n1404 0.0845
R13799 VSS.n1403 VSS.n1402 0.0845
R13800 VSS.n1401 VSS.n1400 0.0845
R13801 VSS.n2075 VSS.n2074 0.0845
R13802 VSS.n2071 VSS.n2070 0.0845
R13803 VSS.n2069 VSS.n2068 0.0845
R13804 VSS.n2067 VSS.n2066 0.0845
R13805 VSS.n702 VSS.n701 0.0845
R13806 VSS.n1506 VSS.n1505 0.0845
R13807 VSS.n1504 VSS.n1503 0.0845
R13808 VSS.n1502 VSS.n1501 0.0845
R13809 VSS.n1500 VSS.n1499 0.0845
R13810 VSS.n1498 VSS.n1497 0.0845
R13811 VSS.n1496 VSS.n1495 0.0845
R13812 VSS.n1494 VSS.n1493 0.0845
R13813 VSS.n1487 VSS.n1486 0.0845
R13814 VSS.n1531 VSS.n1530 0.0845
R13815 VSS.n1529 VSS.n1528 0.0845
R13816 VSS.n449 VSS.n448 0.0845
R13817 VSS.n2083 VSS.n2082 0.0845
R13818 VSS.n2135 VSS.n2134 0.0845
R13819 VSS.n1915 VSS.n1914 0.08375
R13820 VSS.n2055 VSS.n2054 0.08375
R13821 VSS.n838 VSS.n837 0.083
R13822 VSS.n2250 VSS.n2249 0.0815
R13823 VSS.n2253 VSS.n2252 0.0815
R13824 VSS.n1145 VSS.n1144 0.0815
R13825 VSS.n1625 VSS.n1624 0.0815
R13826 VSS.n1621 VSS.n1620 0.0815
R13827 VSS.n1178 VSS.n1177 0.0815
R13828 VSS.n1208 VSS.n1207 0.0815
R13829 VSS.n1268 VSS.n1267 0.0815
R13830 VSS.n1298 VSS.n1297 0.0815
R13831 VSS.n1328 VSS.n1327 0.0815
R13832 VSS.n1966 VSS.n1965 0.0815
R13833 VSS.n1399 VSS.n1398 0.0815
R13834 VSS.n1429 VSS.n1428 0.0815
R13835 VSS.n1508 VSS.n1507 0.0815
R13836 VSS.n1551 VSS.n1541 0.0815
R13837 VSS.n2195 VSS.n2194 0.0815
R13838 VSS.n451 VSS.n450 0.0815
R13839 VSS.n1450 VSS.n1449 0.0815
R13840 VSS.n2530 VSS.n2529 0.0815
R13841 VSS.n2543 VSS.n12 0.0815
R13842 VSS.n2216 VSS.n373 0.0815
R13843 VSS.n2123 VSS.n2122 0.08
R13844 VSS.n965 VSS.n964 0.0785
R13845 VSS.n949 VSS.n948 0.077
R13846 VSS.n1886 VSS.n891 0.077
R13847 VSS.n2406 VSS.n84 0.0755
R13848 VSS.n2404 VSS.n86 0.0755
R13849 VSS.n1738 VSS.n1737 0.07475
R13850 VSS.n1748 VSS.n1747 0.074
R13851 VSS.n2348 VSS.n2347 0.0725
R13852 VSS.n2351 VSS.n2350 0.0725
R13853 VSS.n1082 VSS.n1081 0.0725
R13854 VSS.n1689 VSS.n1688 0.0725
R13855 VSS.n1735 VSS.n1734 0.0725
R13856 VSS.n2174 VSS.n407 0.0725
R13857 VSS.n510 VSS.n405 0.0725
R13858 VSS.n2462 VSS.n56 0.066875
R13859 VSS.n109 VSS.n103 0.066875
R13860 VSS.n138 VSS.n132 0.066875
R13861 VSS.n167 VSS.n161 0.066875
R13862 VSS.n196 VSS.n190 0.066875
R13863 VSS.n225 VSS.n219 0.066875
R13864 VSS.n254 VSS.n248 0.066875
R13865 VSS.n316 VSS.n310 0.066875
R13866 VSS.n1993 VSS.n1990 0.06575
R13867 VSS.n2060 VSS.n2059 0.06575
R13868 VSS.n2465 VSS.n52 0.065132
R13869 VSS.n2469 VSS.n52 0.065132
R13870 VSS.n2470 VSS.n2469 0.065132
R13871 VSS.n2471 VSS.n2470 0.065132
R13872 VSS.n2471 VSS.n49 0.065132
R13873 VSS.n2490 VSS.n50 0.065132
R13874 VSS.n106 VSS.n105 0.064625
R13875 VSS.n135 VSS.n134 0.064625
R13876 VSS.n164 VSS.n163 0.064625
R13877 VSS.n193 VSS.n192 0.064625
R13878 VSS.n222 VSS.n221 0.064625
R13879 VSS.n251 VSS.n250 0.064625
R13880 VSS.n313 VSS.n312 0.064625
R13881 VSS.n2459 VSS.n2458 0.064625
R13882 VSS.n841 VSS.n840 0.062
R13883 VSS.n1042 VSS.n1041 0.0605
R13884 VSS.n1040 VSS.n1039 0.0605
R13885 VSS.n1038 VSS.n1037 0.0605
R13886 VSS.n1036 VSS.n1035 0.0605
R13887 VSS.n1034 VSS.n1033 0.0605
R13888 VSS.n1032 VSS.n1031 0.0605
R13889 VSS.n1030 VSS.n1029 0.0605
R13890 VSS.n996 VSS.n995 0.0605
R13891 VSS.n994 VSS.n993 0.0605
R13892 VSS.n2022 VSS.n2021 0.0605
R13893 VSS.n683 VSS.n682 0.0605
R13894 VSS.n2198 VSS.n387 0.0605
R13895 VSS.n585 VSS.n584 0.0605
R13896 VSS.n1432 VSS.n633 0.0605
R13897 VSS.n2150 VSS.n2149 0.0605
R13898 VSS.n1918 VSS.n1917 0.05975
R13899 VSS.n2184 VSS.n2183 0.05975
R13900 VSS.n1970 VSS.n1969 0.05825
R13901 VSS.n2491 VSS.n49 0.058184
R13902 VSS.n2475 VSS.n50 0.0575377
R13903 VSS.n2041 VSS.n2040 0.0575
R13904 VSS.n356 VSS.n355 0.0565682
R13905 VSS.n346 VSS.n54 0.0565682
R13906 VSS.n2552 VSS.n3 0.0555987
R13907 VSS.n1056 VSS.n1055 0.0545
R13908 VSS.n1730 VSS.n1729 0.0545
R13909 VSS.n1778 VSS.n1777 0.0545
R13910 VSS.n1850 VSS.n893 0.0545
R13911 VSS.n1902 VSS.n1901 0.0545
R13912 VSS.n886 VSS.n885 0.0545
R13913 VSS.n1921 VSS.n1920 0.0545
R13914 VSS.n2048 VSS.n2047 0.0545
R13915 VSS.n740 VSS.n739 0.0545
R13916 VSS.n1528 VSS.n1527 0.0545
R13917 VSS.n2084 VSS.n2083 0.0545
R13918 VSS.n107 VSS.n104 0.0539756
R13919 VSS.n136 VSS.n133 0.0539756
R13920 VSS.n165 VSS.n162 0.0539756
R13921 VSS.n194 VSS.n191 0.0539756
R13922 VSS.n223 VSS.n220 0.0539756
R13923 VSS.n252 VSS.n249 0.0539756
R13924 VSS.n314 VSS.n311 0.0539756
R13925 VSS.n2460 VSS.n57 0.0539756
R13926 VSS.n1983 VSS.n1982 0.05375
R13927 VSS.n2465 VSS.n2464 0.0530135
R13928 VSS.n2312 VSS.n2311 0.0515
R13929 VSS.n1114 VSS.n1113 0.0515
R13930 VSS.n1657 VSS.n1656 0.0515
R13931 VSS.n1713 VSS.n1015 0.0515
R13932 VSS.n1728 VSS.n1727 0.0515
R13933 VSS.n1590 VSS.n1589 0.0515
R13934 VSS.n1742 VSS.n1741 0.0515
R13935 VSS.n1002 VSS.n1001 0.0515
R13936 VSS.n1799 VSS.n1798 0.0515
R13937 VSS.n1803 VSS.n1802 0.0515
R13938 VSS.n1237 VSS.n1236 0.0515
R13939 VSS.n1942 VSS.n1941 0.0515
R13940 VSS.n813 VSS.n812 0.0515
R13941 VSS.n1946 VSS.n1945 0.0515
R13942 VSS.n1369 VSS.n1368 0.0515
R13943 VSS.n2077 VSS.n2076 0.0515
R13944 VSS.n667 VSS.n666 0.0515
R13945 VSS.n572 VSS.n571 0.0515
R13946 VSS.n2200 VSS.n385 0.0515
R13947 VSS.n2486 VSS.n2485 0.0492971
R13948 VSS.n1010 VSS.n1009 0.04925
R13949 VSS.n2044 VSS.n2043 0.0485
R13950 VSS.n1475 VSS.n1474 0.0485
R13951 VSS.n444 VSS.n443 0.0485
R13952 VSS.n354 VSS.n353 0.0483276
R13953 VSS.n1482 VSS.n1481 0.04775
R13954 VSS.n2011 VSS.n2010 0.0455
R13955 VSS.n2032 VSS.n2031 0.0455
R13956 VSS.n2053 VSS.n2052 0.0455
R13957 VSS.n1524 VSS.n1523 0.0455
R13958 VSS.n348 VSS.n347 0.0434802
R13959 VSS.n1737 VSS.n1736 0.04325
R13960 VSS.n108 VSS.n102 0.0426622
R13961 VSS.n137 VSS.n131 0.0426622
R13962 VSS.n166 VSS.n160 0.0426622
R13963 VSS.n195 VSS.n189 0.0426622
R13964 VSS.n224 VSS.n218 0.0426622
R13965 VSS.n253 VSS.n247 0.0426622
R13966 VSS.n315 VSS.n309 0.0426622
R13967 VSS.n2461 VSS.n55 0.0426622
R13968 VSS.n2480 VSS.n2479 0.0425108
R13969 VSS.n294 VSS.n293 0.041125
R13970 VSS.n1835 VSS.n1834 0.041
R13971 VSS.n295 VSS.n258 0.040375
R13972 VSS.n295 VSS.n294 0.039875
R13973 VSS.n2049 VSS.n706 0.0395
R13974 VSS.n2508 VSS.n2498 0.0393636
R13975 VSS.n1553 VSS.n1552 0.0378333
R13976 VSS.n1554 VSS.n1553 0.0378333
R13977 VSS.n1555 VSS.n1554 0.0378333
R13978 VSS.n1556 VSS.n1555 0.0378333
R13979 VSS.n1557 VSS.n1556 0.0378333
R13980 VSS.n1558 VSS.n1557 0.0378333
R13981 VSS.n1559 VSS.n1558 0.0378333
R13982 VSS.n1560 VSS.n1559 0.0378333
R13983 VSS.n1561 VSS.n1560 0.0378333
R13984 VSS.n1562 VSS.n1561 0.0378333
R13985 VSS.n1563 VSS.n1562 0.0378333
R13986 VSS.n1563 VSS.n1147 0.0378333
R13987 VSS.n1147 VSS.n1146 0.0378333
R13988 VSS.n1146 VSS.n95 0.0378333
R13989 VSS.n358 VSS.n95 0.0378333
R13990 VSS.n1734 VSS.n1733 0.03725
R13991 VSS.n2484 VSS.n2483 0.0363707
R13992 VSS.n1749 VSS.n1748 0.03575
R13993 VSS.n2531 VSS.n0 0.0357078
R13994 VSS.n352 VSS.n342 0.0354013
R13995 VSS.n957 VSS.n956 0.03425
R13996 VSS.n734 VSS.n733 0.03425
R13997 VSS.n690 VSS.n689 0.03425
R13998 VSS.n2312 VSS.n93 0.0335
R13999 VSS.n1115 VSS.n1114 0.0335
R14000 VSS.n1656 VSS.n1654 0.0335
R14001 VSS.n1591 VSS.n1590 0.0335
R14002 VSS.n1799 VSS.n911 0.0335
R14003 VSS.n1802 VSS.n909 0.0335
R14004 VSS.n1866 VSS.n1865 0.0335
R14005 VSS.n1238 VSS.n1237 0.0335
R14006 VSS.n1895 VSS.n1894 0.0335
R14007 VSS.n1942 VSS.n780 0.0335
R14008 VSS.n1945 VSS.n778 0.0335
R14009 VSS.n1979 VSS.n1978 0.0335
R14010 VSS.n2077 VSS.n635 0.0335
R14011 VSS.n1013 VSS.n1012 0.03275
R14012 VSS.n1365 VSS.n1364 0.0305
R14013 VSS.n349 VSS.n342 0.0302307
R14014 VSS.n2483 VSS.n2482 0.0292612
R14015 VSS.n1746 VSS.n1745 0.02825
R14016 VSS.n1913 VSS.n1912 0.0275
R14017 VSS.n850 VSS.n849 0.0275
R14018 VSS.n692 VSS.n691 0.0275
R14019 VSS.n1974 VSS.n1973 0.02675
R14020 VSS.n737 VSS.n736 0.02675
R14021 VSS.n2165 VSS.n2164 0.02675
R14022 VSS.n2087 VSS.n2086 0.02675
R14023 VSS.n45 VSS.n22 0.02534
R14024 VSS.n1743 VSS.n1742 0.0245
R14025 VSS.n1831 VSS.n1830 0.0245
R14026 VSS.n1864 VSS.n1863 0.0245
R14027 VSS.n2026 VSS.n2025 0.0245
R14028 VSS.n1908 VSS.n1907 0.02375
R14029 VSS.n2482 VSS.n2480 0.0231212
R14030 VSS.n349 VSS.n348 0.0221517
R14031 VSS.n298 VSS.n297 0.0213379
R14032 VSS.n297 VSS.n258 0.0207356
R14033 VSS.n1875 VSS.n1874 0.01925
R14034 VSS.n2173 VSS.n2172 0.01925
R14035 VSS.n2107 VSS.n2106 0.01925
R14036 VSS.n2144 VSS.n2143 0.01925
R14037 VSS.n844 VSS.n843 0.01775
R14038 VSS.n353 VSS.n352 0.0173043
R14039 VSS.n2485 VSS.n2484 0.0163348
R14040 VSS.n357 VSS.n97 0.0158846
R14041 VSS.n351 VSS.n97 0.0158846
R14042 VSS.n351 VSS.n350 0.0158846
R14043 VSS.n350 VSS.n343 0.0158846
R14044 VSS.n343 VSS.n53 0.0158846
R14045 VSS.n2466 VSS.n53 0.0158846
R14046 VSS.n2467 VSS.n2466 0.0158846
R14047 VSS.n2468 VSS.n2467 0.0158846
R14048 VSS.n2468 VSS.n51 0.0158846
R14049 VSS.n2472 VSS.n51 0.0158846
R14050 VSS.n2473 VSS.n2472 0.0158846
R14051 VSS.n2489 VSS.n2473 0.0158846
R14052 VSS.n2489 VSS.n2488 0.0158846
R14053 VSS.n2488 VSS.n2487 0.0158846
R14054 VSS.n2487 VSS.n2474 0.0158846
R14055 VSS.n2481 VSS.n2474 0.0158846
R14056 VSS.n2481 VSS.n1 0.0158846
R14057 VSS.n2553 VSS.n1 0.0158846
R14058 VSS.n1356 VSS.n1355 0.01325
R14059 VSS.n1489 VSS.n1488 0.01325
R14060 VSS.n2464 VSS.n54 0.0126185
R14061 VSS.n1768 VSS.n1767 0.0125
R14062 VSS.n1908 VSS.n852 0.0125
R14063 VSS.n2186 VSS.n2185 0.01175
R14064 VSS.n2102 VSS.n2101 0.01175
R14065 VSS.n745 VSS.n744 0.011
R14066 VSS.n2479 VSS.n3 0.0100332
R14067 VSS.n355 VSS.n354 0.00906373
R14068 VSS.n347 VSS.n346 0.00906373
R14069 VSS.n1757 VSS.n1756 0.00875
R14070 VSS.n2486 VSS.n2475 0.00809425
R14071 VSS.n2491 VSS.n2490 0.00744794
R14072 VSS.n1349 VSS.n1348 0.0035
R14073 VSS.n2095 VSS.n2094 0.0035
R14074 VSS.n820 VSS.n819 0.00275
R14075 VSS.n674 VSS.n673 0.00275
R14076 VSS.n565 VSS.n564 0.00275
R14077 VSS.n108 VSS.n107 0.00131081
R14078 VSS.n110 VSS.n102 0.00131081
R14079 VSS.n137 VSS.n136 0.00131081
R14080 VSS.n139 VSS.n131 0.00131081
R14081 VSS.n166 VSS.n165 0.00131081
R14082 VSS.n168 VSS.n160 0.00131081
R14083 VSS.n195 VSS.n194 0.00131081
R14084 VSS.n197 VSS.n189 0.00131081
R14085 VSS.n224 VSS.n223 0.00131081
R14086 VSS.n226 VSS.n218 0.00131081
R14087 VSS.n253 VSS.n252 0.00131081
R14088 VSS.n255 VSS.n247 0.00131081
R14089 VSS.n315 VSS.n314 0.00131081
R14090 VSS.n317 VSS.n309 0.00131081
R14091 VSS.n2461 VSS.n2460 0.00131081
R14092 VSS.n2463 VSS.n55 0.00131081
R14093 a_11023_n6840.n2 a_11023_n6840.t26 56.019
R14094 a_11023_n6840.n1 a_11023_n6840.t36 55.9719
R14095 a_11023_n6840.n1 a_11023_n6840.t25 55.9719
R14096 a_11023_n6840.n1 a_11023_n6840.t21 55.9719
R14097 a_11023_n6840.n1 a_11023_n6840.t33 55.9719
R14098 a_11023_n6840.n1 a_11023_n6840.t23 55.9719
R14099 a_11023_n6840.n1 a_11023_n6840.t38 55.9719
R14100 a_11023_n6840.n1 a_11023_n6840.t29 55.9719
R14101 a_11023_n6840.n1 a_11023_n6840.t24 55.9719
R14102 a_11023_n6840.n1 a_11023_n6840.t20 55.9719
R14103 a_11023_n6840.n2 a_11023_n6840.t35 55.9719
R14104 a_11023_n6840.n2 a_11023_n6840.t31 55.9719
R14105 a_11023_n6840.n2 a_11023_n6840.t28 55.9719
R14106 a_11023_n6840.n2 a_11023_n6840.t37 55.9719
R14107 a_11023_n6840.n2 a_11023_n6840.t32 55.9719
R14108 a_11023_n6840.n2 a_11023_n6840.t22 55.9719
R14109 a_11023_n6840.n2 a_11023_n6840.t34 55.9719
R14110 a_11023_n6840.n2 a_11023_n6840.t30 55.9719
R14111 a_11023_n6840.n2 a_11023_n6840.t39 55.9719
R14112 a_11023_n6840.n1 a_11023_n6840.n0 0.14323
R14113 a_11023_n6840.n3 a_11023_n6840.t16 3.87048
R14114 a_11023_n6840.n3 a_11023_n6840.t10 3.68704
R14115 a_11023_n6840.n4 a_11023_n6840.t4 3.68704
R14116 a_11023_n6840.n5 a_11023_n6840.t2 3.68704
R14117 a_11023_n6840.n6 a_11023_n6840.t17 3.68704
R14118 a_11023_n6840.t14 a_11023_n6840.n11 3.53694
R14119 a_11023_n6840.n8 a_11023_n6840.t5 3.37808
R14120 a_11023_n6840.n9 a_11023_n6840.t11 3.37808
R14121 a_11023_n6840.n10 a_11023_n6840.t13 3.37808
R14122 a_11023_n6840.n11 a_11023_n6840.t18 3.37808
R14123 a_11023_n6840.t5 a_11023_n6840.t9 0.6505
R14124 a_11023_n6840.t11 a_11023_n6840.t15 0.6505
R14125 a_11023_n6840.t13 a_11023_n6840.t19 0.6505
R14126 a_11023_n6840.t18 a_11023_n6840.t8 0.6505
R14127 a_11023_n6840.t3 a_11023_n6840.t14 0.6505
R14128 a_11023_n6840.t16 a_11023_n6840.t6 0.5855
R14129 a_11023_n6840.t10 a_11023_n6840.t0 0.5855
R14130 a_11023_n6840.t4 a_11023_n6840.t12 0.5855
R14131 a_11023_n6840.t2 a_11023_n6840.t7 0.5855
R14132 a_11023_n6840.t17 a_11023_n6840.t1 0.5855
R14133 a_11023_n6840.n7 a_11023_n6840.n6 0.41138
R14134 a_11023_n6840.n8 a_11023_n6840.n7 0.373278
R14135 a_11023_n6840.n4 a_11023_n6840.n3 0.183939
R14136 a_11023_n6840.n5 a_11023_n6840.n4 0.183939
R14137 a_11023_n6840.n6 a_11023_n6840.n5 0.183939
R14138 a_11023_n6840.n11 a_11023_n6840.n10 0.159616
R14139 a_11023_n6840.n10 a_11023_n6840.n9 0.159616
R14140 a_11023_n6840.n9 a_11023_n6840.n8 0.159616
R14141 a_11023_n6840.n1 a_11023_n6840.t27 56.3117
R14142 a_11023_n6840.n7 a_11023_n6840.n0 2.08751
R14143 a_11023_n6840.n0 a_11023_n6840.n2 2.43655
R14144 a_13501_n6460.n0 a_13501_n6460.t5 15.8618
R14145 a_13501_n6460.n0 a_13501_n6460.t3 15.8393
R14146 a_13501_n6460.n0 a_13501_n6460.t7 15.7537
R14147 a_13501_n6460.n0 a_13501_n6460.t9 15.7496
R14148 a_13501_n6460.n0 a_13501_n6460.t1 14.963
R14149 a_13501_n6460.n0 a_13501_n6460.t4 14.9583
R14150 a_13501_n6460.n0 a_13501_n6460.t2 14.9559
R14151 a_13501_n6460.n0 a_13501_n6460.t0 14.9547
R14152 a_13501_n6460.n0 a_13501_n6460.t10 14.8524
R14153 a_13501_n6460.n0 a_13501_n6460.t11 14.7096
R14154 a_13501_n6460.t6 a_13501_n6460.n0 14.7035
R14155 a_13501_n6460.n0 a_13501_n6460.t8 14.7035
R14156 a_11087_n7460.n10 a_11087_n7460.t30 12.6085
R14157 a_11087_n7460.n2 a_11087_n7460.n0 10.553
R14158 a_11087_n7460.n10 a_11087_n7460.n9 10.4369
R14159 a_11087_n7460.n12 a_11087_n7460.n11 10.4369
R14160 a_11087_n7460.n14 a_11087_n7460.n13 10.4308
R14161 a_11087_n7460.n16 a_11087_n7460.n15 10.4308
R14162 a_11087_n7460.n18 a_11087_n7460.n17 10.4308
R14163 a_11087_n7460.n2 a_11087_n7460.n1 10.4156
R14164 a_11087_n7460.n6 a_11087_n7460.n5 10.4129
R14165 a_11087_n7460.n8 a_11087_n7460.n7 10.4121
R14166 a_11087_n7460.n4 a_11087_n7460.n3 10.4121
R14167 a_11087_n7460.n28 a_11087_n7460.n27 10.357
R14168 a_11087_n7460.n21 a_11087_n7460.n20 10.2004
R14169 a_11087_n7460.n25 a_11087_n7460.n24 10.2004
R14170 a_11087_n7460.n23 a_11087_n7460.n22 10.198
R14171 a_11087_n7460.n27 a_11087_n7460.n26 10.1921
R14172 a_11087_n7460.n21 a_11087_n7460.n19 0.773592
R14173 a_11087_n7460.n20 a_11087_n7460.t25 0.6505
R14174 a_11087_n7460.n20 a_11087_n7460.t21 0.6505
R14175 a_11087_n7460.n22 a_11087_n7460.t22 0.6505
R14176 a_11087_n7460.n22 a_11087_n7460.t28 0.6505
R14177 a_11087_n7460.n24 a_11087_n7460.t20 0.6505
R14178 a_11087_n7460.n24 a_11087_n7460.t27 0.6505
R14179 a_11087_n7460.n26 a_11087_n7460.t26 0.6505
R14180 a_11087_n7460.n26 a_11087_n7460.t23 0.6505
R14181 a_11087_n7460.n28 a_11087_n7460.t24 0.6505
R14182 a_11087_n7460.t29 a_11087_n7460.n28 0.6505
R14183 a_11087_n7460.n7 a_11087_n7460.t2 0.5855
R14184 a_11087_n7460.n7 a_11087_n7460.t6 0.5855
R14185 a_11087_n7460.n5 a_11087_n7460.t5 0.5855
R14186 a_11087_n7460.n5 a_11087_n7460.t9 0.5855
R14187 a_11087_n7460.n3 a_11087_n7460.t7 0.5855
R14188 a_11087_n7460.n3 a_11087_n7460.t0 0.5855
R14189 a_11087_n7460.n1 a_11087_n7460.t1 0.5855
R14190 a_11087_n7460.n1 a_11087_n7460.t4 0.5855
R14191 a_11087_n7460.n0 a_11087_n7460.t3 0.5855
R14192 a_11087_n7460.n0 a_11087_n7460.t8 0.5855
R14193 a_11087_n7460.n9 a_11087_n7460.t12 0.5855
R14194 a_11087_n7460.n9 a_11087_n7460.t18 0.5855
R14195 a_11087_n7460.n11 a_11087_n7460.t17 0.5855
R14196 a_11087_n7460.n11 a_11087_n7460.t15 0.5855
R14197 a_11087_n7460.n13 a_11087_n7460.t14 0.5855
R14198 a_11087_n7460.n13 a_11087_n7460.t11 0.5855
R14199 a_11087_n7460.n15 a_11087_n7460.t13 0.5855
R14200 a_11087_n7460.n15 a_11087_n7460.t19 0.5855
R14201 a_11087_n7460.n17 a_11087_n7460.t10 0.5855
R14202 a_11087_n7460.n17 a_11087_n7460.t16 0.5855
R14203 a_11087_n7460.n19 a_11087_n7460.n8 0.365893
R14204 a_11087_n7460.n19 a_11087_n7460.n18 0.297718
R14205 a_11087_n7460.n12 a_11087_n7460.n10 0.1615
R14206 a_11087_n7460.n23 a_11087_n7460.n21 0.161
R14207 a_11087_n7460.n18 a_11087_n7460.n16 0.1605
R14208 a_11087_n7460.n16 a_11087_n7460.n14 0.1605
R14209 a_11087_n7460.n27 a_11087_n7460.n25 0.1605
R14210 a_11087_n7460.n25 a_11087_n7460.n23 0.1605
R14211 a_11087_n7460.n14 a_11087_n7460.n12 0.1585
R14212 a_11087_n7460.n8 a_11087_n7460.n6 0.139126
R14213 a_11087_n7460.n4 a_11087_n7460.n2 0.136566
R14214 a_11087_n7460.n6 a_11087_n7460.n4 0.13486
R14215 a_21772_n8292.n5 a_21772_n8292.t23 15.8415
R14216 a_21772_n8292.n6 a_21772_n8292.t13 15.8415
R14217 a_21772_n8292.n7 a_21772_n8292.t11 15.8415
R14218 a_21772_n8292.n8 a_21772_n8292.t14 15.8415
R14219 a_21772_n8292.n9 a_21772_n8292.t16 15.8415
R14220 a_21772_n8292.n10 a_21772_n8292.t19 15.8415
R14221 a_21772_n8292.n4 a_21772_n8292.t18 15.8415
R14222 a_21772_n8292.n11 a_21772_n8292.t20 15.8415
R14223 a_21772_n8292.n5 a_21772_n8292.t17 13.4447
R14224 a_21772_n8292.n6 a_21772_n8292.t21 13.4447
R14225 a_21772_n8292.n7 a_21772_n8292.t22 13.4447
R14226 a_21772_n8292.n8 a_21772_n8292.t8 13.4447
R14227 a_21772_n8292.n9 a_21772_n8292.t10 13.4447
R14228 a_21772_n8292.n10 a_21772_n8292.t9 13.4447
R14229 a_21772_n8292.n4 a_21772_n8292.t12 13.4447
R14230 a_21772_n8292.n11 a_21772_n8292.t15 13.4447
R14231 a_21772_n8292.n6 a_21772_n8292.n5 10.5449
R14232 a_21772_n8292.n7 a_21772_n8292.n6 10.5449
R14233 a_21772_n8292.n8 a_21772_n8292.n7 10.5449
R14234 a_21772_n8292.n9 a_21772_n8292.n8 10.5449
R14235 a_21772_n8292.n10 a_21772_n8292.n9 10.5449
R14236 a_21772_n8292.n11 a_21772_n8292.n4 10.5449
R14237 a_21772_n8292.n11 a_21772_n8292.n10 10.5449
R14238 a_21772_n8292.n0 a_21772_n8292.n3 7.22489
R14239 a_21772_n8292.n0 a_21772_n8292.n2 6.36702
R14240 a_21772_n8292.n12 a_21772_n8292.n0 3.56115
R14241 a_21772_n8292.n0 a_21772_n8292.n1 2.68463
R14242 a_21772_n8292.n0 a_21772_n8292.n11 2.37183
R14243 a_21772_n8292.n1 a_21772_n8292.t4 2.06607
R14244 a_21772_n8292.t7 a_21772_n8292.n12 2.06607
R14245 a_21772_n8292.n2 a_21772_n8292.t2 1.99806
R14246 a_21772_n8292.n2 a_21772_n8292.t3 1.99806
R14247 a_21772_n8292.n3 a_21772_n8292.t0 1.99806
R14248 a_21772_n8292.n3 a_21772_n8292.t1 1.99806
R14249 a_21772_n8292.n1 a_21772_n8292.t5 1.4923
R14250 a_21772_n8292.n12 a_21772_n8292.t6 1.4923
R14251 a_13623_n17552.n0 a_13623_n17552.t42 56.1018
R14252 a_13623_n17552.n2 a_13623_n17552.t44 56.0719
R14253 a_13623_n17552.n0 a_13623_n17552.t38 56.0141
R14254 a_13623_n17552.n0 a_13623_n17552.t23 55.9719
R14255 a_13623_n17552.n0 a_13623_n17552.t35 55.9719
R14256 a_13623_n17552.n0 a_13623_n17552.t45 55.9719
R14257 a_13623_n17552.n0 a_13623_n17552.t28 55.9719
R14258 a_13623_n17552.n0 a_13623_n17552.t20 55.9719
R14259 a_13623_n17552.n0 a_13623_n17552.t30 55.9719
R14260 a_13623_n17552.n0 a_13623_n17552.t41 55.9719
R14261 a_13623_n17552.n0 a_13623_n17552.t22 55.9719
R14262 a_13623_n17552.n0 a_13623_n17552.t34 55.9719
R14263 a_13623_n17552.n0 a_13623_n17552.t18 55.9719
R14264 a_13623_n17552.n0 a_13623_n17552.t32 55.9719
R14265 a_13623_n17552.n0 a_13623_n17552.t39 55.9719
R14266 a_13623_n17552.n0 a_13623_n17552.t25 55.9719
R14267 a_13623_n17552.n0 a_13623_n17552.t16 55.9719
R14268 a_13623_n17552.n0 a_13623_n17552.t26 55.9719
R14269 a_13623_n17552.n0 a_13623_n17552.t37 55.9719
R14270 a_13623_n17552.n0 a_13623_n17552.t17 55.9719
R14271 a_13623_n17552.n0 a_13623_n17552.t31 55.9719
R14272 a_13623_n17552.n2 a_13623_n17552.t27 55.9719
R14273 a_13623_n17552.n2 a_13623_n17552.t36 55.9719
R14274 a_13623_n17552.n2 a_13623_n17552.t29 55.9719
R14275 a_13623_n17552.n2 a_13623_n17552.t40 55.9719
R14276 a_13623_n17552.n2 a_13623_n17552.t21 55.9719
R14277 a_13623_n17552.n2 a_13623_n17552.t33 55.9719
R14278 a_13623_n17552.n4 a_13623_n17552.t43 55.9719
R14279 a_13623_n17552.n4 a_13623_n17552.t24 55.9719
R14280 a_13623_n17552.n4 a_13623_n17552.t19 55.9719
R14281 a_13623_n17552.n3 a_13623_n17552.n0 38.9545
R14282 a_13623_n17552.n1 a_13623_n17552.n8 6.90733
R14283 a_13623_n17552.n1 a_13623_n17552.n10 6.89497
R14284 a_13623_n17552.n1 a_13623_n17552.n9 6.3768
R14285 a_13623_n17552.n1 a_13623_n17552.n7 6.3768
R14286 a_13623_n17552.n1 a_13623_n17552.n6 3.21104
R14287 a_13623_n17552.n3 a_13623_n17552.n11 2.83209
R14288 a_13623_n17552.n1 a_13623_n17552.n5 2.7042
R14289 a_13623_n17552.n12 a_13623_n17552.n1 2.7042
R14290 a_13623_n17552.n6 a_13623_n17552.t11 2.06607
R14291 a_13623_n17552.n5 a_13623_n17552.t12 2.06607
R14292 a_13623_n17552.n11 a_13623_n17552.t8 2.06607
R14293 a_13623_n17552.t15 a_13623_n17552.n12 2.06607
R14294 a_13623_n17552.n9 a_13623_n17552.t6 1.99806
R14295 a_13623_n17552.n9 a_13623_n17552.t5 1.99806
R14296 a_13623_n17552.n10 a_13623_n17552.t4 1.99806
R14297 a_13623_n17552.n10 a_13623_n17552.t3 1.99806
R14298 a_13623_n17552.n8 a_13623_n17552.t1 1.99806
R14299 a_13623_n17552.n8 a_13623_n17552.t2 1.99806
R14300 a_13623_n17552.n7 a_13623_n17552.t7 1.99806
R14301 a_13623_n17552.n7 a_13623_n17552.t0 1.99806
R14302 a_13623_n17552.n6 a_13623_n17552.t9 1.4923
R14303 a_13623_n17552.n5 a_13623_n17552.t10 1.4923
R14304 a_13623_n17552.n11 a_13623_n17552.t14 1.4923
R14305 a_13623_n17552.n12 a_13623_n17552.t13 1.4923
R14306 a_13623_n17552.n1 a_13623_n17552.n3 1.23036
R14307 a_13623_n17552.n0 a_13623_n17552.n4 1.21455
R14308 a_13623_n17552.n4 a_13623_n17552.n2 0.8005
R14309 a_11023_n14874.n2 a_11023_n14874.t38 56.019
R14310 a_11023_n14874.n1 a_11023_n14874.t26 55.9719
R14311 a_11023_n14874.n1 a_11023_n14874.t34 55.9719
R14312 a_11023_n14874.n1 a_11023_n14874.t21 55.9719
R14313 a_11023_n14874.n1 a_11023_n14874.t36 55.9719
R14314 a_11023_n14874.n1 a_11023_n14874.t23 55.9719
R14315 a_11023_n14874.n1 a_11023_n14874.t30 55.9719
R14316 a_11023_n14874.n1 a_11023_n14874.t39 55.9719
R14317 a_11023_n14874.n1 a_11023_n14874.t25 55.9719
R14318 a_11023_n14874.n1 a_11023_n14874.t31 55.9719
R14319 a_11023_n14874.n2 a_11023_n14874.t27 55.9719
R14320 a_11023_n14874.n2 a_11023_n14874.t33 55.9719
R14321 a_11023_n14874.n2 a_11023_n14874.t20 55.9719
R14322 a_11023_n14874.n2 a_11023_n14874.t28 55.9719
R14323 a_11023_n14874.n2 a_11023_n14874.t35 55.9719
R14324 a_11023_n14874.n2 a_11023_n14874.t22 55.9719
R14325 a_11023_n14874.n2 a_11023_n14874.t37 55.9719
R14326 a_11023_n14874.n2 a_11023_n14874.t24 55.9719
R14327 a_11023_n14874.n2 a_11023_n14874.t32 55.9719
R14328 a_11023_n14874.n1 a_11023_n14874.n0 0.14323
R14329 a_11023_n14874.n4 a_11023_n14874.t15 3.87048
R14330 a_11023_n14874.n4 a_11023_n14874.t0 3.68704
R14331 a_11023_n14874.n5 a_11023_n14874.t6 3.68704
R14332 a_11023_n14874.n6 a_11023_n14874.t2 3.68704
R14333 a_11023_n14874.n7 a_11023_n14874.t8 3.68704
R14334 a_11023_n14874.n3 a_11023_n14874.t13 3.53719
R14335 a_11023_n14874.n9 a_11023_n14874.t5 3.37808
R14336 a_11023_n14874.n10 a_11023_n14874.t19 3.37808
R14337 a_11023_n14874.n3 a_11023_n14874.t17 3.37808
R14338 a_11023_n14874.t9 a_11023_n14874.n11 3.37783
R14339 a_11023_n14874.t5 a_11023_n14874.t18 0.6505
R14340 a_11023_n14874.t19 a_11023_n14874.t14 0.6505
R14341 a_11023_n14874.t17 a_11023_n14874.t10 0.6505
R14342 a_11023_n14874.t13 a_11023_n14874.t4 0.6505
R14343 a_11023_n14874.t3 a_11023_n14874.t9 0.6505
R14344 a_11023_n14874.t15 a_11023_n14874.t7 0.5855
R14345 a_11023_n14874.t0 a_11023_n14874.t12 0.5855
R14346 a_11023_n14874.t6 a_11023_n14874.t11 0.5855
R14347 a_11023_n14874.t2 a_11023_n14874.t16 0.5855
R14348 a_11023_n14874.t8 a_11023_n14874.t1 0.5855
R14349 a_11023_n14874.n8 a_11023_n14874.n7 0.41138
R14350 a_11023_n14874.n9 a_11023_n14874.n8 0.373278
R14351 a_11023_n14874.n5 a_11023_n14874.n4 0.183939
R14352 a_11023_n14874.n6 a_11023_n14874.n5 0.183939
R14353 a_11023_n14874.n7 a_11023_n14874.n6 0.183939
R14354 a_11023_n14874.n11 a_11023_n14874.n3 0.159616
R14355 a_11023_n14874.n11 a_11023_n14874.n10 0.159616
R14356 a_11023_n14874.n10 a_11023_n14874.n9 0.159616
R14357 a_11023_n14874.n1 a_11023_n14874.t29 56.3117
R14358 a_11023_n14874.n8 a_11023_n14874.n0 2.08751
R14359 a_11023_n14874.n0 a_11023_n14874.n2 2.43655
R14360 a_11087_n15494.n26 a_11087_n15494.t33 14.158
R14361 a_11087_n15494.n27 a_11087_n15494.n26 14.0623
R14362 a_11087_n15494.n12 a_11087_n15494.n10 10.553
R14363 a_11087_n15494.n29 a_11087_n15494.n28 10.4369
R14364 a_11087_n15494.n31 a_11087_n15494.n30 10.4369
R14365 a_11087_n15494.n25 a_11087_n15494.n24 10.4308
R14366 a_11087_n15494.n23 a_11087_n15494.n22 10.4308
R14367 a_11087_n15494.n21 a_11087_n15494.n20 10.4308
R14368 a_11087_n15494.n12 a_11087_n15494.n11 10.4156
R14369 a_11087_n15494.n16 a_11087_n15494.n15 10.4129
R14370 a_11087_n15494.n18 a_11087_n15494.n17 10.4121
R14371 a_11087_n15494.n14 a_11087_n15494.n13 10.4121
R14372 a_11087_n15494.n3 a_11087_n15494.n1 10.357
R14373 a_11087_n15494.n9 a_11087_n15494.n8 10.2004
R14374 a_11087_n15494.n5 a_11087_n15494.n4 10.2004
R14375 a_11087_n15494.n7 a_11087_n15494.n6 10.198
R14376 a_11087_n15494.n3 a_11087_n15494.n2 10.1921
R14377 a_11087_n15494.n29 a_11087_n15494.n27 2.57417
R14378 a_11087_n15494.n26 a_11087_n15494.t32 1.07268
R14379 a_11087_n15494.n19 a_11087_n15494.n9 0.773592
R14380 a_11087_n15494.n8 a_11087_n15494.t12 0.6505
R14381 a_11087_n15494.n8 a_11087_n15494.t16 0.6505
R14382 a_11087_n15494.n6 a_11087_n15494.t11 0.6505
R14383 a_11087_n15494.n6 a_11087_n15494.t19 0.6505
R14384 a_11087_n15494.n4 a_11087_n15494.t14 0.6505
R14385 a_11087_n15494.n4 a_11087_n15494.t18 0.6505
R14386 a_11087_n15494.n2 a_11087_n15494.t17 0.6505
R14387 a_11087_n15494.n2 a_11087_n15494.t10 0.6505
R14388 a_11087_n15494.n1 a_11087_n15494.t15 0.6505
R14389 a_11087_n15494.n1 a_11087_n15494.t13 0.6505
R14390 a_11087_n15494.n28 a_11087_n15494.t26 0.5855
R14391 a_11087_n15494.n28 a_11087_n15494.t20 0.5855
R14392 a_11087_n15494.n24 a_11087_n15494.t22 0.5855
R14393 a_11087_n15494.n24 a_11087_n15494.t25 0.5855
R14394 a_11087_n15494.n22 a_11087_n15494.t21 0.5855
R14395 a_11087_n15494.n22 a_11087_n15494.t28 0.5855
R14396 a_11087_n15494.n20 a_11087_n15494.t24 0.5855
R14397 a_11087_n15494.n20 a_11087_n15494.t27 0.5855
R14398 a_11087_n15494.n17 a_11087_n15494.t6 0.5855
R14399 a_11087_n15494.n17 a_11087_n15494.t2 0.5855
R14400 a_11087_n15494.n15 a_11087_n15494.t7 0.5855
R14401 a_11087_n15494.n15 a_11087_n15494.t9 0.5855
R14402 a_11087_n15494.n13 a_11087_n15494.t4 0.5855
R14403 a_11087_n15494.n13 a_11087_n15494.t0 0.5855
R14404 a_11087_n15494.n11 a_11087_n15494.t1 0.5855
R14405 a_11087_n15494.n11 a_11087_n15494.t8 0.5855
R14406 a_11087_n15494.n10 a_11087_n15494.t3 0.5855
R14407 a_11087_n15494.n10 a_11087_n15494.t5 0.5855
R14408 a_11087_n15494.t29 a_11087_n15494.n31 0.5855
R14409 a_11087_n15494.n31 a_11087_n15494.t23 0.5855
R14410 a_11087_n15494.n19 a_11087_n15494.n18 0.366893
R14411 a_11087_n15494.n0 a_11087_n15494.t30 10.6208
R14412 a_11087_n15494.n21 a_11087_n15494.n19 0.297718
R14413 a_11087_n15494.n30 a_11087_n15494.n29 0.1615
R14414 a_11087_n15494.n9 a_11087_n15494.n7 0.161
R14415 a_11087_n15494.n5 a_11087_n15494.n3 0.1605
R14416 a_11087_n15494.n7 a_11087_n15494.n5 0.1605
R14417 a_11087_n15494.n23 a_11087_n15494.n21 0.1605
R14418 a_11087_n15494.n25 a_11087_n15494.n23 0.1605
R14419 a_11087_n15494.n30 a_11087_n15494.n25 0.1585
R14420 a_11087_n15494.n18 a_11087_n15494.n16 0.139126
R14421 a_11087_n15494.n14 a_11087_n15494.n12 0.136566
R14422 a_11087_n15494.n16 a_11087_n15494.n14 0.13486
R14423 a_11087_n15494.n0 a_11087_n15494.t31 1.02798
R14424 a_11087_n15494.n27 a_11087_n15494.n0 11.4264
R14425 a_28721_n9076.n4 a_28721_n9076.t5 22.1195
R14426 a_28721_n9076.n3 a_28721_n9076.n2 21.6805
R14427 a_28721_n9076.n3 a_28721_n9076.n1 19.9261
R14428 a_28721_n9076.n5 a_28721_n9076.t2 19.5645
R14429 a_28721_n9076.n2 a_28721_n9076.t7 19.4185
R14430 a_28721_n9076.n1 a_28721_n9076.t6 18.6885
R14431 a_28721_n9076.n5 a_28721_n9076.t8 18.4938
R14432 a_28721_n9076.t1 a_28721_n9076.n0 17.7305
R14433 a_28721_n9076.n1 a_28721_n9076.t3 11.9603
R14434 a_28721_n9076.n2 a_28721_n9076.t4 11.6683
R14435 a_28721_n9076.n0 a_28721_n9076.n3 10.0805
R14436 a_28721_n9076.t1 a_28721_n9076.t0 9.85539
R14437 a_28721_n9076.n4 a_28721_n9076.t9 9.02817
R14438 a_28721_n9076.n0 a_28721_n9076.n5 8.51318
R14439 a_28721_n9076.n0 a_28721_n9076.n4 8.35407
R14440 a_26440_n5940.n2 a_26440_n5940.t7 15.7685
R14441 a_26440_n5940.n3 a_26440_n5940.t16 15.7685
R14442 a_26440_n5940.n4 a_26440_n5940.t9 15.7685
R14443 a_26440_n5940.n5 a_26440_n5940.t5 15.7685
R14444 a_26440_n5940.n6 a_26440_n5940.t13 15.7685
R14445 a_26440_n5940.n7 a_26440_n5940.t6 15.7685
R14446 a_26440_n5940.n1 a_26440_n5940.t11 15.7685
R14447 a_26440_n5940.n0 a_26440_n5940.t14 15.7685
R14448 a_26440_n5940.n0 a_26440_n5940.t3 12.3783
R14449 a_26440_n5940.n2 a_26440_n5940.t10 11.6197
R14450 a_26440_n5940.n3 a_26440_n5940.t12 11.6197
R14451 a_26440_n5940.n4 a_26440_n5940.t15 11.6197
R14452 a_26440_n5940.n5 a_26440_n5940.t17 11.6197
R14453 a_26440_n5940.n6 a_26440_n5940.t19 11.6197
R14454 a_26440_n5940.n7 a_26440_n5940.t18 11.6197
R14455 a_26440_n5940.n1 a_26440_n5940.t8 11.6197
R14456 a_26440_n5940.n0 a_26440_n5940.t4 11.6197
R14457 a_26440_n5940.n3 a_26440_n5940.n2 10.5449
R14458 a_26440_n5940.n4 a_26440_n5940.n3 10.5449
R14459 a_26440_n5940.n5 a_26440_n5940.n4 10.5449
R14460 a_26440_n5940.n6 a_26440_n5940.n5 10.5449
R14461 a_26440_n5940.n7 a_26440_n5940.n6 10.5449
R14462 a_26440_n5940.n0 a_26440_n5940.n1 10.5449
R14463 a_26440_n5940.n0 a_26440_n5940.t2 10.4819
R14464 a_26440_n5940.n0 a_26440_n5940.t1 9.32628
R14465 a_26440_n5940.t0 a_26440_n5940.n0 8.44976
R14466 a_26440_n5940.n0 a_26440_n5940.n7 8.41578
R14467 a_21692_n5468.n21 a_21692_n5468.n20 18.7205
R14468 a_21692_n5468.n21 a_21692_n5468.n5 17.7988
R14469 a_21692_n5468.n12 a_21692_n5468.n11 17.5073
R14470 a_21692_n5468.n9 a_21692_n5468.n7 14.0423
R14471 a_21692_n5468.n11 a_21692_n5468.t19 13.615
R14472 a_21692_n5468.n6 a_21692_n5468.t26 13.615
R14473 a_21692_n5468.n8 a_21692_n5468.t16 13.615
R14474 a_21692_n5468.n19 a_21692_n5468.t24 13.5542
R14475 a_21692_n5468.n17 a_21692_n5468.t18 13.5542
R14476 a_21692_n5468.n15 a_21692_n5468.t22 13.5542
R14477 a_21692_n5468.n7 a_21692_n5468.t27 13.5542
R14478 a_21692_n5468.n13 a_21692_n5468.t21 13.1892
R14479 a_21692_n5468.n5 a_21692_n5468.t28 13.1892
R14480 a_21692_n5468.n10 a_21692_n5468.n6 13.0073
R14481 a_21692_n5468.n13 a_21692_n5468.t17 12.8485
R14482 a_21692_n5468.n5 a_21692_n5468.t20 12.8485
R14483 a_21692_n5468.n9 a_21692_n5468.n8 12.8273
R14484 a_21692_n5468.n14 a_21692_n5468.n13 12.6238
R14485 a_21692_n5468.n20 a_21692_n5468.n19 12.6189
R14486 a_21692_n5468.n16 a_21692_n5468.n15 12.6189
R14487 a_21692_n5468.n18 a_21692_n5468.n17 12.5147
R14488 a_21692_n5468.n19 a_21692_n5468.t33 12.4105
R14489 a_21692_n5468.n17 a_21692_n5468.t25 12.4105
R14490 a_21692_n5468.n15 a_21692_n5468.t30 12.4105
R14491 a_21692_n5468.n7 a_21692_n5468.t31 12.4105
R14492 a_21692_n5468.n11 a_21692_n5468.t23 12.3375
R14493 a_21692_n5468.n6 a_21692_n5468.t29 12.3375
R14494 a_21692_n5468.n8 a_21692_n5468.t32 12.3375
R14495 a_21692_n5468.n12 a_21692_n5468.n10 10.6205
R14496 a_21692_n5468.n14 a_21692_n5468.n12 9.43866
R14497 a_21692_n5468.n2 a_21692_n5468.n25 7.13263
R14498 a_21692_n5468.n1 a_21692_n5468.n23 7.13263
R14499 a_21692_n5468.n2 a_21692_n5468.n24 6.43746
R14500 a_21692_n5468.n1 a_21692_n5468.n22 6.43746
R14501 a_21692_n5468.n18 a_21692_n5468.n16 5.1305
R14502 a_21692_n5468.n0 a_21692_n5468.n21 4.6805
R14503 a_21692_n5468.n16 a_21692_n5468.n14 4.1405
R14504 a_21692_n5468.n25 a_21692_n5468.t6 3.8098
R14505 a_21692_n5468.n25 a_21692_n5468.t7 3.8098
R14506 a_21692_n5468.n24 a_21692_n5468.t1 3.8098
R14507 a_21692_n5468.n24 a_21692_n5468.t0 3.8098
R14508 a_21692_n5468.n22 a_21692_n5468.t2 3.8098
R14509 a_21692_n5468.n22 a_21692_n5468.t3 3.8098
R14510 a_21692_n5468.n23 a_21692_n5468.t4 3.8098
R14511 a_21692_n5468.n23 a_21692_n5468.t5 3.8098
R14512 a_21692_n5468.n0 a_21692_n5468.n26 3.34593
R14513 a_21692_n5468.n0 a_21692_n5468.n4 2.80031
R14514 a_21692_n5468.n0 a_21692_n5468.n3 2.71593
R14515 a_21692_n5468.n27 a_21692_n5468.n0 2.71593
R14516 a_21692_n5468.n20 a_21692_n5468.n18 2.6555
R14517 a_21692_n5468.n10 a_21692_n5468.n9 2.1155
R14518 a_21692_n5468.n3 a_21692_n5468.t14 2.06607
R14519 a_21692_n5468.n3 a_21692_n5468.t10 2.06607
R14520 a_21692_n5468.n4 a_21692_n5468.t11 2.06607
R14521 a_21692_n5468.n4 a_21692_n5468.t9 2.06607
R14522 a_21692_n5468.n26 a_21692_n5468.t8 2.06607
R14523 a_21692_n5468.n26 a_21692_n5468.t13 2.06607
R14524 a_21692_n5468.t15 a_21692_n5468.n27 2.06607
R14525 a_21692_n5468.n27 a_21692_n5468.t12 2.06607
R14526 a_21692_n5468.n0 a_21692_n5468.n1 1.3428
R14527 a_21692_n5468.n1 a_21692_n5468.n2 0.577741
R14528 a_11023_n17552.n21 a_11023_n17552.t25 56.0276
R14529 a_11023_n17552.n10 a_11023_n17552.t34 56.019
R14530 a_11023_n17552.n12 a_11023_n17552.t22 55.9719
R14531 a_11023_n17552.n6 a_11023_n17552.t30 55.9719
R14532 a_11023_n17552.n14 a_11023_n17552.t37 55.9719
R14533 a_11023_n17552.n5 a_11023_n17552.t32 55.9719
R14534 a_11023_n17552.n16 a_11023_n17552.t39 55.9719
R14535 a_11023_n17552.n4 a_11023_n17552.t26 55.9719
R14536 a_11023_n17552.n17 a_11023_n17552.t35 55.9719
R14537 a_11023_n17552.n2 a_11023_n17552.t21 55.9719
R14538 a_11023_n17552.n22 a_11023_n17552.t27 55.9719
R14539 a_11023_n17552.n10 a_11023_n17552.t23 55.9719
R14540 a_11023_n17552.n10 a_11023_n17552.t29 55.9719
R14541 a_11023_n17552.n9 a_11023_n17552.t36 55.9719
R14542 a_11023_n17552.n9 a_11023_n17552.t24 55.9719
R14543 a_11023_n17552.n7 a_11023_n17552.t31 55.9719
R14544 a_11023_n17552.n7 a_11023_n17552.t38 55.9719
R14545 a_11023_n17552.n8 a_11023_n17552.t33 55.9719
R14546 a_11023_n17552.n8 a_11023_n17552.t20 55.9719
R14547 a_11023_n17552.n27 a_11023_n17552.t28 55.9719
R14548 a_11023_n17552.n12 a_11023_n17552.n11 0.0590857
R14549 a_11023_n17552.n24 a_11023_n17552.n23 4.5005
R14550 a_11023_n17552.n25 a_11023_n17552.n2 4.5005
R14551 a_11023_n17552.n17 a_11023_n17552.n26 4.5005
R14552 a_11023_n17552.n3 a_11023_n17552.n0 4.5005
R14553 a_11023_n17552.n1 a_11023_n17552.n4 4.5005
R14554 a_11023_n17552.n16 a_11023_n17552.n15 4.5005
R14555 a_11023_n17552.n33 a_11023_n17552.n32 4.5005
R14556 a_11023_n17552.n31 a_11023_n17552.n5 4.5005
R14557 a_11023_n17552.n14 a_11023_n17552.n13 4.5005
R14558 a_11023_n17552.n30 a_11023_n17552.n29 4.5005
R14559 a_11023_n17552.n28 a_11023_n17552.n6 4.5005
R14560 a_11023_n17552.n39 a_11023_n17552.n38 3.87048
R14561 a_11023_n17552.n39 a_11023_n17552.n37 3.68704
R14562 a_11023_n17552.n40 a_11023_n17552.n36 3.68704
R14563 a_11023_n17552.n41 a_11023_n17552.n35 3.68704
R14564 a_11023_n17552.n42 a_11023_n17552.n34 3.68704
R14565 a_11023_n17552.n20 a_11023_n17552.n18 3.53719
R14566 a_11023_n17552.n45 a_11023_n17552.n44 3.37808
R14567 a_11023_n17552.n47 a_11023_n17552.n46 3.37808
R14568 a_11023_n17552.n20 a_11023_n17552.n19 3.37808
R14569 a_11023_n17552.n49 a_11023_n17552.n48 3.37783
R14570 a_11023_n17552.n43 a_11023_n17552.n1 1.89107
R14571 a_11023_n17552.n24 a_11023_n17552.n21 1.15666
R14572 a_11023_n17552.n44 a_11023_n17552.t17 0.6505
R14573 a_11023_n17552.n44 a_11023_n17552.t11 0.6505
R14574 a_11023_n17552.n46 a_11023_n17552.t10 0.6505
R14575 a_11023_n17552.n46 a_11023_n17552.t13 0.6505
R14576 a_11023_n17552.n19 a_11023_n17552.t12 0.6505
R14577 a_11023_n17552.n19 a_11023_n17552.t15 0.6505
R14578 a_11023_n17552.n18 a_11023_n17552.t14 0.6505
R14579 a_11023_n17552.n18 a_11023_n17552.t18 0.6505
R14580 a_11023_n17552.t19 a_11023_n17552.n49 0.6505
R14581 a_11023_n17552.n49 a_11023_n17552.t16 0.6505
R14582 a_11023_n17552.n38 a_11023_n17552.t4 0.5855
R14583 a_11023_n17552.n38 a_11023_n17552.t8 0.5855
R14584 a_11023_n17552.n37 a_11023_n17552.t2 0.5855
R14585 a_11023_n17552.n37 a_11023_n17552.t5 0.5855
R14586 a_11023_n17552.n36 a_11023_n17552.t9 0.5855
R14587 a_11023_n17552.n36 a_11023_n17552.t6 0.5855
R14588 a_11023_n17552.n35 a_11023_n17552.t0 0.5855
R14589 a_11023_n17552.n35 a_11023_n17552.t3 0.5855
R14590 a_11023_n17552.n34 a_11023_n17552.t7 0.5855
R14591 a_11023_n17552.n34 a_11023_n17552.t1 0.5855
R14592 a_11023_n17552.n43 a_11023_n17552.n42 0.41138
R14593 a_11023_n17552.n45 a_11023_n17552.n43 0.373278
R14594 a_11023_n17552.n40 a_11023_n17552.n39 0.183939
R14595 a_11023_n17552.n41 a_11023_n17552.n40 0.183939
R14596 a_11023_n17552.n42 a_11023_n17552.n41 0.183939
R14597 a_11023_n17552.n48 a_11023_n17552.n20 0.159616
R14598 a_11023_n17552.n48 a_11023_n17552.n47 0.159616
R14599 a_11023_n17552.n47 a_11023_n17552.n45 0.159616
R14600 a_11023_n17552.n22 a_11023_n17552.n21 0.121859
R14601 a_11023_n17552.n23 a_11023_n17552.n22 0.11975
R14602 a_11023_n17552.n17 a_11023_n17552.n2 0.11975
R14603 a_11023_n17552.n4 a_11023_n17552.n16 0.11975
R14604 a_11023_n17552.n5 a_11023_n17552.n14 0.11975
R14605 a_11023_n17552.n6 a_11023_n17552.n12 0.11975
R14606 a_11023_n17552.n25 a_11023_n17552.n24 0.11975
R14607 a_11023_n17552.n26 a_11023_n17552.n25 0.11975
R14608 a_11023_n17552.n26 a_11023_n17552.n0 0.11975
R14609 a_11023_n17552.n1 a_11023_n17552.n15 0.11975
R14610 a_11023_n17552.n32 a_11023_n17552.n15 0.11975
R14611 a_11023_n17552.n32 a_11023_n17552.n31 0.11975
R14612 a_11023_n17552.n31 a_11023_n17552.n13 0.11975
R14613 a_11023_n17552.n29 a_11023_n17552.n13 0.11975
R14614 a_11023_n17552.n29 a_11023_n17552.n28 0.11975
R14615 a_11023_n17552.n28 a_11023_n17552.n11 2.37025
R14616 a_11023_n17552.n3 a_11023_n17552.n17 0.11975
R14617 a_11023_n17552.n16 a_11023_n17552.n33 0.11975
R14618 a_11023_n17552.n14 a_11023_n17552.n30 0.11975
R14619 a_11023_n17552.n11 a_11023_n17552.n27 1.35571
R14620 a_11023_n17552.n30 a_11023_n17552.n6 0.11975
R14621 a_11023_n17552.n33 a_11023_n17552.n5 0.11975
R14622 a_11023_n17552.n4 a_11023_n17552.n3 0.11975
R14623 a_11023_n17552.n23 a_11023_n17552.n2 0.11975
R14624 a_11023_n17552.n1 a_11023_n17552.n0 0.11975
R14625 a_11023_n17552.n9 a_11023_n17552.n10 0.0946176
R14626 a_11023_n17552.n7 a_11023_n17552.n9 0.0946176
R14627 a_11023_n17552.n8 a_11023_n17552.n7 0.0946176
R14628 a_11023_n17552.n27 a_11023_n17552.n8 0.0946176
R14629 a_11087_n18172.n25 a_11087_n18172.n22 17.2039
R14630 a_11087_n18172.n13 a_11087_n18172.n11 10.553
R14631 a_11087_n18172.n27 a_11087_n18172.n26 10.4369
R14632 a_11087_n18172.n29 a_11087_n18172.n28 10.4369
R14633 a_11087_n18172.n31 a_11087_n18172.n30 10.4308
R14634 a_11087_n18172.n33 a_11087_n18172.n32 10.4308
R14635 a_11087_n18172.n35 a_11087_n18172.n34 10.4308
R14636 a_11087_n18172.n13 a_11087_n18172.n12 10.4156
R14637 a_11087_n18172.n17 a_11087_n18172.n16 10.4129
R14638 a_11087_n18172.n19 a_11087_n18172.n18 10.4121
R14639 a_11087_n18172.n15 a_11087_n18172.n14 10.4121
R14640 a_11087_n18172.n4 a_11087_n18172.n2 10.357
R14641 a_11087_n18172.n10 a_11087_n18172.n9 10.2004
R14642 a_11087_n18172.n6 a_11087_n18172.n5 10.2004
R14643 a_11087_n18172.n8 a_11087_n18172.n7 10.198
R14644 a_11087_n18172.n4 a_11087_n18172.n3 10.1921
R14645 a_11087_n18172.n1 a_11087_n18172.n23 6.22845
R14646 a_11087_n18172.n0 a_11087_n18172.n21 6.22852
R14647 a_11087_n18172.n25 a_11087_n18172.n24 5.00122
R14648 a_11087_n18172.n27 a_11087_n18172.n25 2.09842
R14649 a_11087_n18172.n22 a_11087_n18172.t36 1.23128
R14650 a_11087_n18172.n23 a_11087_n18172.t34 1.21988
R14651 a_11087_n18172.n24 a_11087_n18172.t31 1.21875
R14652 a_11087_n18172.n21 a_11087_n18172.t33 1.2147
R14653 a_11087_n18172.n20 a_11087_n18172.n10 0.773592
R14654 a_11087_n18172.n9 a_11087_n18172.t14 0.6505
R14655 a_11087_n18172.n9 a_11087_n18172.t18 0.6505
R14656 a_11087_n18172.n7 a_11087_n18172.t13 0.6505
R14657 a_11087_n18172.n7 a_11087_n18172.t11 0.6505
R14658 a_11087_n18172.n5 a_11087_n18172.t16 0.6505
R14659 a_11087_n18172.n5 a_11087_n18172.t10 0.6505
R14660 a_11087_n18172.n3 a_11087_n18172.t19 0.6505
R14661 a_11087_n18172.n3 a_11087_n18172.t12 0.6505
R14662 a_11087_n18172.n2 a_11087_n18172.t17 0.6505
R14663 a_11087_n18172.n2 a_11087_n18172.t15 0.6505
R14664 a_11087_n18172.n26 a_11087_n18172.t28 0.5855
R14665 a_11087_n18172.n26 a_11087_n18172.t22 0.5855
R14666 a_11087_n18172.n28 a_11087_n18172.t21 0.5855
R14667 a_11087_n18172.n28 a_11087_n18172.t25 0.5855
R14668 a_11087_n18172.n30 a_11087_n18172.t24 0.5855
R14669 a_11087_n18172.n30 a_11087_n18172.t27 0.5855
R14670 a_11087_n18172.n32 a_11087_n18172.t23 0.5855
R14671 a_11087_n18172.n32 a_11087_n18172.t20 0.5855
R14672 a_11087_n18172.n18 a_11087_n18172.t6 0.5855
R14673 a_11087_n18172.n18 a_11087_n18172.t0 0.5855
R14674 a_11087_n18172.n16 a_11087_n18172.t5 0.5855
R14675 a_11087_n18172.n16 a_11087_n18172.t3 0.5855
R14676 a_11087_n18172.n14 a_11087_n18172.t8 0.5855
R14677 a_11087_n18172.n14 a_11087_n18172.t2 0.5855
R14678 a_11087_n18172.n12 a_11087_n18172.t1 0.5855
R14679 a_11087_n18172.n12 a_11087_n18172.t4 0.5855
R14680 a_11087_n18172.n11 a_11087_n18172.t9 0.5855
R14681 a_11087_n18172.n11 a_11087_n18172.t7 0.5855
R14682 a_11087_n18172.n35 a_11087_n18172.t26 0.5855
R14683 a_11087_n18172.t29 a_11087_n18172.n35 0.5855
R14684 a_11087_n18172.n20 a_11087_n18172.n19 0.366893
R14685 a_11087_n18172.n21 a_11087_n18172.t35 7.26093
R14686 a_11087_n18172.n1 a_11087_n18172.t30 1.02798
R14687 a_11087_n18172.n23 a_11087_n18172.t37 7.24134
R14688 a_11087_n18172.n34 a_11087_n18172.n20 0.297718
R14689 a_11087_n18172.n29 a_11087_n18172.n27 0.1615
R14690 a_11087_n18172.n10 a_11087_n18172.n8 0.161
R14691 a_11087_n18172.n6 a_11087_n18172.n4 0.1605
R14692 a_11087_n18172.n8 a_11087_n18172.n6 0.1605
R14693 a_11087_n18172.n34 a_11087_n18172.n33 0.1605
R14694 a_11087_n18172.n33 a_11087_n18172.n31 0.1605
R14695 a_11087_n18172.n31 a_11087_n18172.n29 0.1585
R14696 a_11087_n18172.n19 a_11087_n18172.n17 0.139126
R14697 a_11087_n18172.n15 a_11087_n18172.n13 0.136566
R14698 a_11087_n18172.n17 a_11087_n18172.n15 0.13486
R14699 a_11087_n18172.n22 a_11087_n18172.n0 6.22741
R14700 a_11087_n18172.n24 a_11087_n18172.n1 6.22829
R14701 a_11087_n18172.n0 a_11087_n18172.t32 1.03316
R14702 a_26388_n17606.t1 a_26388_n17606.n9 33.8855
R14703 a_26388_n17606.n1 a_26388_n17606.n2 23.1275
R14704 a_26388_n17606.n9 a_26388_n17606.n7 21.7355
R14705 a_26388_n17606.n1 a_26388_n17606.n5 19.8455
R14706 a_26388_n17606.n2 a_26388_n17606.t7 19.5645
R14707 a_26388_n17606.n8 a_26388_n17606.t8 17.4475
R14708 a_26388_n17606.n4 a_26388_n17606.t10 17.192
R14709 a_26388_n17606.n2 a_26388_n17606.t5 17.1312
R14710 a_26388_n17606.n5 a_26388_n17606.n3 15.3005
R14711 a_26388_n17606.n9 a_26388_n17606.n8 12.8393
R14712 a_26388_n17606.n8 a_26388_n17606.t11 12.7755
R14713 a_26388_n17606.n4 a_26388_n17606.t3 12.3497
R14714 a_26388_n17606.n7 a_26388_n17606.n1 10.6366
R14715 a_26388_n17606.t1 a_26388_n17606.t0 9.70112
R14716 a_26388_n17606.n5 a_26388_n17606.n4 8.5545
R14717 a_26388_n17606.n0 a_26388_n17606.t9 6.71423
R14718 a_26388_n17606.n3 a_26388_n17606.t13 6.71423
R14719 a_26388_n17606.n6 a_26388_n17606.t2 6.3005
R14720 a_26388_n17606.n6 a_26388_n17606.t12 5.6196
R14721 a_26388_n17606.n0 a_26388_n17606.t6 5.20587
R14722 a_26388_n17606.n3 a_26388_n17606.t4 5.20587
R14723 a_26388_n17606.n7 a_26388_n17606.n6 4.71811
R14724 a_26388_n17606.n1 a_26388_n17606.n0 4.6805
R14725 a_10778_2852.n0 a_10778_2852.t26 55.9719
R14726 a_10778_2852.n0 a_10778_2852.t21 55.9719
R14727 a_10778_2852.n0 a_10778_2852.t18 55.9719
R14728 a_10778_2852.n0 a_10778_2852.t32 55.9719
R14729 a_10778_2852.n0 a_10778_2852.t19 55.9719
R14730 a_10778_2852.n0 a_10778_2852.t34 55.9719
R14731 a_10778_2852.n0 a_10778_2852.t30 55.9719
R14732 a_10778_2852.n0 a_10778_2852.t27 55.9719
R14733 a_10778_2852.n0 a_10778_2852.t24 55.9719
R14734 a_10778_2852.n0 a_10778_2852.t22 55.9719
R14735 a_10778_2852.n0 a_10778_2852.t20 55.9719
R14736 a_10778_2852.n0 a_10778_2852.t15 55.9719
R14737 a_10778_2852.n0 a_10778_2852.t31 55.9719
R14738 a_10778_2852.n0 a_10778_2852.t28 55.9719
R14739 a_10778_2852.n0 a_10778_2852.t33 55.9719
R14740 a_10778_2852.n0 a_10778_2852.t29 55.9719
R14741 a_10778_2852.n0 a_10778_2852.t25 55.9719
R14742 a_10778_2852.n0 a_10778_2852.t23 55.9719
R14743 a_10778_2852.n0 a_10778_2852.t17 55.9719
R14744 a_10778_2852.n0 a_10778_2852.t16 55.9719
R14745 a_10778_2852.n2 a_10778_2852.t11 9.42441
R14746 a_10778_2852.n1 a_10778_2852.t10 9.42441
R14747 a_10778_2852.n1 a_10778_2852.t12 9.42441
R14748 a_10778_2852.n1 a_10778_2852.t13 9.42441
R14749 a_10778_2852.n1 a_10778_2852.t14 9.42441
R14750 a_10778_2852.n2 a_10778_2852.n0 8.42934
R14751 a_10778_2852.n2 a_10778_2852.t5 8.15873
R14752 a_10778_2852.n1 a_10778_2852.t4 8.15873
R14753 a_10778_2852.n1 a_10778_2852.t9 8.15873
R14754 a_10778_2852.n1 a_10778_2852.t2 8.15873
R14755 a_10778_2852.n1 a_10778_2852.t0 8.15873
R14756 a_10778_2852.n3 a_10778_2852.t6 8.14399
R14757 a_10778_2852.t1 a_10778_2852.n3 7.93973
R14758 a_10778_2852.n3 a_10778_2852.t8 7.93973
R14759 a_10778_2852.n3 a_10778_2852.t7 7.93973
R14760 a_10778_2852.n3 a_10778_2852.t3 7.93973
R14761 a_10778_2852.n2 a_10778_2852.n1 1.32239
R14762 a_10778_2852.n3 a_10778_2852.n2 0.941067
R14763 a_10712_4516.n9 a_10712_4516.n7 59.2654
R14764 a_10712_4516.n1 a_10712_4516.t46 55.9719
R14765 a_10712_4516.n4 a_10712_4516.t41 55.9719
R14766 a_10712_4516.n4 a_10712_4516.t40 55.9719
R14767 a_10712_4516.n3 a_10712_4516.t42 55.9719
R14768 a_10712_4516.n3 a_10712_4516.t36 55.9719
R14769 a_10712_4516.n2 a_10712_4516.t33 55.9719
R14770 a_10712_4516.n2 a_10712_4516.t52 55.9719
R14771 a_10712_4516.n0 a_10712_4516.t50 55.9719
R14772 a_10712_4516.n0 a_10712_4516.t45 55.9719
R14773 a_10712_4516.n1 a_10712_4516.t48 55.9719
R14774 a_10712_4516.n4 a_10712_4516.t34 55.9719
R14775 a_10712_4516.n4 a_10712_4516.t32 55.9719
R14776 a_10712_4516.n3 a_10712_4516.t35 55.9719
R14777 a_10712_4516.n3 a_10712_4516.t53 55.9719
R14778 a_10712_4516.n2 a_10712_4516.t51 55.9719
R14779 a_10712_4516.n2 a_10712_4516.t47 55.9719
R14780 a_10712_4516.n0 a_10712_4516.t44 55.9719
R14781 a_10712_4516.n0 a_10712_4516.t37 55.9719
R14782 a_10712_4516.n1 a_10712_4516.t39 55.9719
R14783 a_10712_4516.n1 a_10712_4516.t38 55.9719
R14784 a_10712_4516.n6 a_10712_4516.t43 19.7105
R14785 a_10712_4516.n6 a_10712_4516.t49 13.3108
R14786 a_10712_4516.n7 a_10712_4516.n6 13.2998
R14787 a_10712_4516.n7 a_10712_4516.n5 12.4205
R14788 a_10712_4516.n28 a_10712_4516.n14 7.35813
R14789 a_10712_4516.n26 a_10712_4516.n15 7.35813
R14790 a_10712_4516.n24 a_10712_4516.n16 7.35813
R14791 a_10712_4516.n22 a_10712_4516.n17 7.35813
R14792 a_10712_4516.n20 a_10712_4516.n18 7.35813
R14793 a_10712_4516.n5 a_10712_4516.t31 6.71423
R14794 a_10712_4516.n28 a_10712_4516.n27 5.90992
R14795 a_10712_4516.n26 a_10712_4516.n25 5.90992
R14796 a_10712_4516.n24 a_10712_4516.n23 5.90992
R14797 a_10712_4516.n22 a_10712_4516.n21 5.90992
R14798 a_10712_4516.n20 a_10712_4516.n19 5.90992
R14799 a_10712_4516.n29 a_10712_4516.n1 5.71583
R14800 a_10712_4516.n31 a_10712_4516.n30 5.69092
R14801 a_10712_4516.n13 a_10712_4516.n12 5.69092
R14802 a_10712_4516.n11 a_10712_4516.n10 5.69092
R14803 a_10712_4516.n9 a_10712_4516.n8 5.69092
R14804 a_10712_4516.n33 a_10712_4516.n32 5.69092
R14805 a_10712_4516.n5 a_10712_4516.t30 5.20587
R14806 a_10712_4516.n30 a_10712_4516.t27 0.6505
R14807 a_10712_4516.n30 a_10712_4516.t24 0.6505
R14808 a_10712_4516.n12 a_10712_4516.t20 0.6505
R14809 a_10712_4516.n12 a_10712_4516.t28 0.6505
R14810 a_10712_4516.n10 a_10712_4516.t23 0.6505
R14811 a_10712_4516.n10 a_10712_4516.t22 0.6505
R14812 a_10712_4516.n8 a_10712_4516.t26 0.6505
R14813 a_10712_4516.n8 a_10712_4516.t25 0.6505
R14814 a_10712_4516.n33 a_10712_4516.t21 0.6505
R14815 a_10712_4516.t29 a_10712_4516.n33 0.6505
R14816 a_10712_4516.n27 a_10712_4516.t19 0.5855
R14817 a_10712_4516.n27 a_10712_4516.t16 0.5855
R14818 a_10712_4516.n14 a_10712_4516.t7 0.5855
R14819 a_10712_4516.n14 a_10712_4516.t0 0.5855
R14820 a_10712_4516.n25 a_10712_4516.t13 0.5855
R14821 a_10712_4516.n25 a_10712_4516.t11 0.5855
R14822 a_10712_4516.n15 a_10712_4516.t3 0.5855
R14823 a_10712_4516.n15 a_10712_4516.t5 0.5855
R14824 a_10712_4516.n23 a_10712_4516.t12 0.5855
R14825 a_10712_4516.n23 a_10712_4516.t10 0.5855
R14826 a_10712_4516.n16 a_10712_4516.t4 0.5855
R14827 a_10712_4516.n16 a_10712_4516.t6 0.5855
R14828 a_10712_4516.n21 a_10712_4516.t15 0.5855
R14829 a_10712_4516.n21 a_10712_4516.t14 0.5855
R14830 a_10712_4516.n17 a_10712_4516.t1 0.5855
R14831 a_10712_4516.n17 a_10712_4516.t2 0.5855
R14832 a_10712_4516.n19 a_10712_4516.t18 0.5855
R14833 a_10712_4516.n19 a_10712_4516.t17 0.5855
R14834 a_10712_4516.n18 a_10712_4516.t8 0.5855
R14835 a_10712_4516.n18 a_10712_4516.t9 0.5855
R14836 a_10712_4516.n31 a_10712_4516.n29 0.39704
R14837 a_10712_4516.n29 a_10712_4516.n28 0.284406
R14838 a_10712_4516.n11 a_10712_4516.n9 0.255367
R14839 a_10712_4516.n13 a_10712_4516.n11 0.255367
R14840 a_10712_4516.n32 a_10712_4516.n13 0.255367
R14841 a_10712_4516.n32 a_10712_4516.n31 0.255367
R14842 a_10712_4516.n22 a_10712_4516.n20 0.223756
R14843 a_10712_4516.n24 a_10712_4516.n22 0.223756
R14844 a_10712_4516.n26 a_10712_4516.n24 0.223756
R14845 a_10712_4516.n28 a_10712_4516.n26 0.223756
R14846 a_10712_4516.n1 a_10712_4516.n0 0.195893
R14847 a_10712_4516.n3 a_10712_4516.n4 0.13023
R14848 a_10712_4516.n2 a_10712_4516.n3 0.13023
R14849 a_10712_4516.n0 a_10712_4516.n2 0.13023
R14850 a_44640_1944.n9 a_44640_1944.t10 15.8415
R14851 a_44640_1944.n3 a_44640_1944.t16 15.8415
R14852 a_44640_1944.n4 a_44640_1944.t17 15.8415
R14853 a_44640_1944.n5 a_44640_1944.t13 15.8415
R14854 a_44640_1944.n6 a_44640_1944.t15 15.8415
R14855 a_44640_1944.n7 a_44640_1944.t11 15.8415
R14856 a_44640_1944.n8 a_44640_1944.t12 15.8415
R14857 a_44640_1944.n10 a_44640_1944.t14 15.8415
R14858 a_44640_1944.n9 a_44640_1944.t18 13.4447
R14859 a_44640_1944.n3 a_44640_1944.t8 13.4447
R14860 a_44640_1944.n4 a_44640_1944.t9 13.4447
R14861 a_44640_1944.n5 a_44640_1944.t21 13.4447
R14862 a_44640_1944.n6 a_44640_1944.t23 13.4447
R14863 a_44640_1944.n7 a_44640_1944.t19 13.4447
R14864 a_44640_1944.n8 a_44640_1944.t20 13.4447
R14865 a_44640_1944.n10 a_44640_1944.t22 13.4447
R14866 a_44640_1944.n4 a_44640_1944.n3 10.5449
R14867 a_44640_1944.n5 a_44640_1944.n4 10.5449
R14868 a_44640_1944.n6 a_44640_1944.n5 10.5449
R14869 a_44640_1944.n7 a_44640_1944.n6 10.5449
R14870 a_44640_1944.n8 a_44640_1944.n7 10.5449
R14871 a_44640_1944.n10 a_44640_1944.n8 10.5449
R14872 a_44640_1944.n10 a_44640_1944.n9 10.5449
R14873 a_44640_1944.n0 a_44640_1944.n2 7.22489
R14874 a_44640_1944.n0 a_44640_1944.n1 6.36702
R14875 a_44640_1944.n0 a_44640_1944.n11 3.56115
R14876 a_44640_1944.n12 a_44640_1944.n0 2.68463
R14877 a_44640_1944.n0 a_44640_1944.n10 2.37181
R14878 a_44640_1944.n11 a_44640_1944.t6 2.06607
R14879 a_44640_1944.n12 a_44640_1944.t4 2.06607
R14880 a_44640_1944.n1 a_44640_1944.t0 1.99806
R14881 a_44640_1944.n1 a_44640_1944.t3 1.99806
R14882 a_44640_1944.n2 a_44640_1944.t2 1.99806
R14883 a_44640_1944.n2 a_44640_1944.t1 1.99806
R14884 a_44640_1944.n11 a_44640_1944.t5 1.4923
R14885 a_44640_1944.t7 a_44640_1944.n12 1.4923
R14886 OUT[5] OUT[5].n14 19.6925
R14887 OUT[5].n3 OUT[5].n2 6.90733
R14888 OUT[5].n3 OUT[5].n1 6.3768
R14889 OUT[5].n12 OUT[5].n0 6.3768
R14890 OUT[5].n14 OUT[5].n13 6.3005
R14891 OUT[5].n9 OUT[5].n8 3.23472
R14892 OUT[5].n6 OUT[5].n5 3.21104
R14893 OUT[5].n9 OUT[5].n7 2.7042
R14894 OUT[5].n6 OUT[5].n4 2.7042
R14895 OUT[5].n7 OUT[5].t12 2.06607
R14896 OUT[5].n8 OUT[5].t9 2.06607
R14897 OUT[5].n5 OUT[5].t15 2.06607
R14898 OUT[5].n4 OUT[5].t14 2.06607
R14899 OUT[5].n13 OUT[5].t1 1.99806
R14900 OUT[5].n13 OUT[5].t5 1.99806
R14901 OUT[5].n2 OUT[5].t7 1.99806
R14902 OUT[5].n2 OUT[5].t6 1.99806
R14903 OUT[5].n1 OUT[5].t2 1.99806
R14904 OUT[5].n1 OUT[5].t0 1.99806
R14905 OUT[5].n0 OUT[5].t4 1.99806
R14906 OUT[5].n0 OUT[5].t3 1.99806
R14907 OUT[5].n7 OUT[5].t10 1.4923
R14908 OUT[5].n8 OUT[5].t8 1.4923
R14909 OUT[5].n5 OUT[5].t11 1.4923
R14910 OUT[5].n4 OUT[5].t13 1.4923
R14911 OUT[5].n14 OUT[5].n12 0.577837
R14912 OUT[5].n11 OUT[5].n3 0.189974
R14913 OUT[5].n10 OUT[5].n6 0.175763
R14914 OUT[5].n10 OUT[5].n9 0.166289
R14915 OUT[5].n12 OUT[5].n11 0.152079
R14916 OUT[5].n11 OUT[5].n10 0.145625
R14917 a_13623_n9518.n0 a_13623_n9518.t36 56.1018
R14918 a_13623_n9518.n0 a_13623_n9518.t23 56.0719
R14919 a_13623_n9518.n0 a_13623_n9518.t18 56.0141
R14920 a_13623_n9518.n0 a_13623_n9518.t29 55.9719
R14921 a_13623_n9518.n0 a_13623_n9518.t14 55.9719
R14922 a_13623_n9518.n0 a_13623_n9518.t37 55.9719
R14923 a_13623_n9518.n0 a_13623_n9518.t20 55.9719
R14924 a_13623_n9518.n0 a_13623_n9518.t9 55.9719
R14925 a_13623_n9518.n0 a_13623_n9518.t33 55.9719
R14926 a_13623_n9518.n0 a_13623_n9518.t16 55.9719
R14927 a_13623_n9518.n0 a_13623_n9518.t12 55.9719
R14928 a_13623_n9518.n0 a_13623_n9518.t24 55.9719
R14929 a_13623_n9518.n0 a_13623_n9518.t27 55.9719
R14930 a_13623_n9518.n0 a_13623_n9518.t11 55.9719
R14931 a_13623_n9518.n0 a_13623_n9518.t19 55.9719
R14932 a_13623_n9518.n0 a_13623_n9518.t32 55.9719
R14933 a_13623_n9518.n0 a_13623_n9518.t25 55.9719
R14934 a_13623_n9518.n0 a_13623_n9518.t34 55.9719
R14935 a_13623_n9518.n0 a_13623_n9518.t17 55.9719
R14936 a_13623_n9518.n0 a_13623_n9518.t26 55.9719
R14937 a_13623_n9518.n0 a_13623_n9518.t10 55.9719
R14938 a_13623_n9518.n0 a_13623_n9518.t35 55.9719
R14939 a_13623_n9518.n0 a_13623_n9518.t15 55.9719
R14940 a_13623_n9518.n0 a_13623_n9518.t8 55.9719
R14941 a_13623_n9518.n0 a_13623_n9518.t21 55.9719
R14942 a_13623_n9518.n0 a_13623_n9518.t30 55.9719
R14943 a_13623_n9518.n0 a_13623_n9518.t13 55.9719
R14944 a_13623_n9518.n0 a_13623_n9518.t22 55.9719
R14945 a_13623_n9518.n0 a_13623_n9518.t31 55.9719
R14946 a_13623_n9518.n0 a_13623_n9518.t28 55.9719
R14947 a_13623_n9518.n1 a_13623_n9518.n0 46.3045
R14948 a_13623_n9518.n1 a_13623_n9518.t5 6.90733
R14949 a_13623_n9518.n1 a_13623_n9518.t0 6.89497
R14950 a_13623_n9518.n1 a_13623_n9518.t7 6.3768
R14951 a_13623_n9518.n1 a_13623_n9518.t1 6.3768
R14952 a_13623_n9518.t2 a_13623_n9518.n1 5.57839
R14953 a_13623_n9518.n1 a_13623_n9518.t3 5.3003
R14954 a_13623_n9518.n1 a_13623_n9518.t6 5.27661
R14955 a_13623_n9518.n1 a_13623_n9518.t4 4.76977
R14956 a_11087_n10138.n4 a_11087_n10138.t20 10.553
R14957 a_11087_n10138.n8 a_11087_n10138.t11 10.4369
R14958 a_11087_n10138.n9 a_11087_n10138.t6 10.4369
R14959 a_11087_n10138.n10 a_11087_n10138.t1 10.4308
R14960 a_11087_n10138.n11 a_11087_n10138.t4 10.4308
R14961 a_11087_n10138.n12 a_11087_n10138.t18 10.4308
R14962 a_11087_n10138.n4 a_11087_n10138.t22 10.4156
R14963 a_11087_n10138.n6 a_11087_n10138.t26 10.4129
R14964 a_11087_n10138.n7 a_11087_n10138.t27 10.4121
R14965 a_11087_n10138.n5 a_11087_n10138.t29 10.4121
R14966 a_11087_n10138.n1 a_11087_n10138.t2 10.357
R14967 a_11087_n10138.n2 a_11087_n10138.t12 10.2004
R14968 a_11087_n10138.t10 a_11087_n10138.n14 10.2004
R14969 a_11087_n10138.n3 a_11087_n10138.t7 10.198
R14970 a_11087_n10138.n1 a_11087_n10138.t17 10.1921
R14971 a_11087_n10138.n14 a_11087_n10138.n13 0.773592
R14972 a_11087_n10138.t7 a_11087_n10138.t15 0.6505
R14973 a_11087_n10138.t12 a_11087_n10138.t16 0.6505
R14974 a_11087_n10138.t17 a_11087_n10138.t3 0.6505
R14975 a_11087_n10138.t2 a_11087_n10138.t14 0.6505
R14976 a_11087_n10138.t0 a_11087_n10138.t10 0.6505
R14977 a_11087_n10138.t27 a_11087_n10138.t21 0.5855
R14978 a_11087_n10138.t26 a_11087_n10138.t24 0.5855
R14979 a_11087_n10138.t29 a_11087_n10138.t23 0.5855
R14980 a_11087_n10138.t22 a_11087_n10138.t25 0.5855
R14981 a_11087_n10138.t20 a_11087_n10138.t28 0.5855
R14982 a_11087_n10138.t11 a_11087_n10138.t5 0.5855
R14983 a_11087_n10138.t6 a_11087_n10138.t19 0.5855
R14984 a_11087_n10138.t1 a_11087_n10138.t13 0.5855
R14985 a_11087_n10138.t4 a_11087_n10138.t8 0.5855
R14986 a_11087_n10138.t18 a_11087_n10138.t9 0.5855
R14987 a_11087_n10138.n13 a_11087_n10138.n7 0.365893
R14988 a_11087_n10138.n0 a_11087_n10138.t30 3.871
R14989 a_11087_n10138.n13 a_11087_n10138.n12 0.297718
R14990 a_11087_n10138.n9 a_11087_n10138.n8 0.1615
R14991 a_11087_n10138.n14 a_11087_n10138.n3 0.161
R14992 a_11087_n10138.n12 a_11087_n10138.n11 0.1605
R14993 a_11087_n10138.n11 a_11087_n10138.n10 0.1605
R14994 a_11087_n10138.n2 a_11087_n10138.n1 0.1605
R14995 a_11087_n10138.n3 a_11087_n10138.n2 0.1605
R14996 a_11087_n10138.n10 a_11087_n10138.n9 0.1585
R14997 a_11087_n10138.n7 a_11087_n10138.n6 0.139126
R14998 a_11087_n10138.n5 a_11087_n10138.n4 0.136566
R14999 a_11087_n10138.n6 a_11087_n10138.n5 0.13486
R15000 a_11087_n10138.n0 a_11087_n10138.t31 1.02798
R15001 a_11087_n10138.n8 a_11087_n10138.n0 17.3038
R15002 a_13501_n9138.n1 a_13501_n9138.t14 15.8618
R15003 a_13501_n9138.n0 a_13501_n9138.t13 15.8393
R15004 a_13501_n9138.n1 a_13501_n9138.t4 15.7537
R15005 a_13501_n9138.n0 a_13501_n9138.t1 15.7496
R15006 a_13501_n9138.n0 a_13501_n9138.n2 14.963
R15007 a_13501_n9138.n9 a_13501_n9138.n1 14.9583
R15008 a_13501_n9138.n1 a_13501_n9138.n5 14.9559
R15009 a_13501_n9138.n1 a_13501_n9138.n6 14.9547
R15010 a_13501_n9138.n0 a_13501_n9138.n3 14.7096
R15011 a_13501_n9138.n1 a_13501_n9138.n7 14.7035
R15012 a_13501_n9138.n1 a_13501_n9138.n8 14.7035
R15013 a_13501_n9138.n1 a_13501_n9138.n4 14.6941
R15014 a_13501_n9138.n4 a_13501_n9138.t7 0.6505
R15015 a_13501_n9138.n4 a_13501_n9138.t0 0.6505
R15016 a_13501_n9138.n7 a_13501_n9138.t8 0.6505
R15017 a_13501_n9138.n7 a_13501_n9138.t3 0.6505
R15018 a_13501_n9138.n8 a_13501_n9138.t2 0.6505
R15019 a_13501_n9138.n8 a_13501_n9138.t5 0.6505
R15020 a_13501_n9138.n3 a_13501_n9138.t6 0.6505
R15021 a_13501_n9138.n3 a_13501_n9138.t9 0.6505
R15022 a_13501_n9138.n5 a_13501_n9138.t17 0.5855
R15023 a_13501_n9138.n5 a_13501_n9138.t10 0.5855
R15024 a_13501_n9138.n6 a_13501_n9138.t16 0.5855
R15025 a_13501_n9138.n6 a_13501_n9138.t19 0.5855
R15026 a_13501_n9138.n2 a_13501_n9138.t11 0.5855
R15027 a_13501_n9138.n2 a_13501_n9138.t15 0.5855
R15028 a_13501_n9138.t18 a_13501_n9138.n9 0.5855
R15029 a_13501_n9138.n9 a_13501_n9138.t12 0.5855
R15030 a_13501_n9138.n1 a_13501_n9138.n0 0.158862
R15031 a_13623_n22908.n0 a_13623_n22908.t25 56.1018
R15032 a_13623_n22908.n0 a_13623_n22908.t27 56.0719
R15033 a_13623_n22908.n0 a_13623_n22908.t21 56.0141
R15034 a_13623_n22908.n0 a_13623_n22908.t36 55.9719
R15035 a_13623_n22908.n0 a_13623_n22908.t18 55.9719
R15036 a_13623_n22908.n0 a_13623_n22908.t28 55.9719
R15037 a_13623_n22908.n0 a_13623_n22908.t11 55.9719
R15038 a_13623_n22908.n0 a_13623_n22908.t33 55.9719
R15039 a_13623_n22908.n0 a_13623_n22908.t13 55.9719
R15040 a_13623_n22908.n0 a_13623_n22908.t24 55.9719
R15041 a_13623_n22908.n0 a_13623_n22908.t35 55.9719
R15042 a_13623_n22908.n0 a_13623_n22908.t17 55.9719
R15043 a_13623_n22908.n0 a_13623_n22908.t31 55.9719
R15044 a_13623_n22908.n0 a_13623_n22908.t15 55.9719
R15045 a_13623_n22908.n0 a_13623_n22908.t22 55.9719
R15046 a_13623_n22908.n0 a_13623_n22908.t8 55.9719
R15047 a_13623_n22908.n0 a_13623_n22908.t29 55.9719
R15048 a_13623_n22908.n0 a_13623_n22908.t9 55.9719
R15049 a_13623_n22908.n0 a_13623_n22908.t20 55.9719
R15050 a_13623_n22908.n0 a_13623_n22908.t30 55.9719
R15051 a_13623_n22908.n0 a_13623_n22908.t14 55.9719
R15052 a_13623_n22908.n0 a_13623_n22908.t10 55.9719
R15053 a_13623_n22908.n0 a_13623_n22908.t19 55.9719
R15054 a_13623_n22908.n0 a_13623_n22908.t12 55.9719
R15055 a_13623_n22908.n0 a_13623_n22908.t23 55.9719
R15056 a_13623_n22908.n0 a_13623_n22908.t34 55.9719
R15057 a_13623_n22908.n0 a_13623_n22908.t16 55.9719
R15058 a_13623_n22908.n0 a_13623_n22908.t26 55.9719
R15059 a_13623_n22908.n0 a_13623_n22908.t37 55.9719
R15060 a_13623_n22908.n0 a_13623_n22908.t32 55.9719
R15061 a_13623_n22908.n1 a_13623_n22908.n0 43.0559
R15062 a_13623_n22908.n1 a_13623_n22908.t4 6.90733
R15063 a_13623_n22908.n1 a_13623_n22908.t7 6.89497
R15064 a_13623_n22908.n1 a_13623_n22908.t6 6.3768
R15065 a_13623_n22908.n1 a_13623_n22908.t5 6.3768
R15066 a_13623_n22908.t0 a_13623_n22908.n1 6.12753
R15067 a_13623_n22908.n1 a_13623_n22908.t3 5.27661
R15068 a_13623_n22908.n1 a_13623_n22908.t1 4.76977
R15069 a_13623_n22908.n1 a_13623_n22908.t2 4.76977
R15070 a_11023_n22908.n21 a_11023_n22908.t38 56.0276
R15071 a_11023_n22908.n10 a_11023_n22908.t27 56.019
R15072 a_11023_n22908.n12 a_11023_n22908.t35 55.9719
R15073 a_11023_n22908.n6 a_11023_n22908.t23 55.9719
R15074 a_11023_n22908.n14 a_11023_n22908.t30 55.9719
R15075 a_11023_n22908.n5 a_11023_n22908.t25 55.9719
R15076 a_11023_n22908.n16 a_11023_n22908.t32 55.9719
R15077 a_11023_n22908.n4 a_11023_n22908.t39 55.9719
R15078 a_11023_n22908.n17 a_11023_n22908.t28 55.9719
R15079 a_11023_n22908.n2 a_11023_n22908.t34 55.9719
R15080 a_11023_n22908.n22 a_11023_n22908.t20 55.9719
R15081 a_11023_n22908.n10 a_11023_n22908.t36 55.9719
R15082 a_11023_n22908.n10 a_11023_n22908.t22 55.9719
R15083 a_11023_n22908.n9 a_11023_n22908.t29 55.9719
R15084 a_11023_n22908.n9 a_11023_n22908.t37 55.9719
R15085 a_11023_n22908.n7 a_11023_n22908.t24 55.9719
R15086 a_11023_n22908.n7 a_11023_n22908.t31 55.9719
R15087 a_11023_n22908.n8 a_11023_n22908.t26 55.9719
R15088 a_11023_n22908.n8 a_11023_n22908.t33 55.9719
R15089 a_11023_n22908.n27 a_11023_n22908.t21 55.9719
R15090 a_11023_n22908.n12 a_11023_n22908.n11 0.0590857
R15091 a_11023_n22908.n24 a_11023_n22908.n23 4.5005
R15092 a_11023_n22908.n25 a_11023_n22908.n2 4.5005
R15093 a_11023_n22908.n17 a_11023_n22908.n26 4.5005
R15094 a_11023_n22908.n3 a_11023_n22908.n0 4.5005
R15095 a_11023_n22908.n1 a_11023_n22908.n4 4.5005
R15096 a_11023_n22908.n16 a_11023_n22908.n15 4.5005
R15097 a_11023_n22908.n33 a_11023_n22908.n32 4.5005
R15098 a_11023_n22908.n31 a_11023_n22908.n5 4.5005
R15099 a_11023_n22908.n14 a_11023_n22908.n13 4.5005
R15100 a_11023_n22908.n30 a_11023_n22908.n29 4.5005
R15101 a_11023_n22908.n28 a_11023_n22908.n6 4.5005
R15102 a_11023_n22908.n39 a_11023_n22908.n38 3.87048
R15103 a_11023_n22908.n39 a_11023_n22908.n37 3.68704
R15104 a_11023_n22908.n40 a_11023_n22908.n36 3.68704
R15105 a_11023_n22908.n41 a_11023_n22908.n35 3.68704
R15106 a_11023_n22908.n42 a_11023_n22908.n34 3.68704
R15107 a_11023_n22908.n20 a_11023_n22908.n18 3.53719
R15108 a_11023_n22908.n45 a_11023_n22908.n44 3.37808
R15109 a_11023_n22908.n47 a_11023_n22908.n46 3.37808
R15110 a_11023_n22908.n20 a_11023_n22908.n19 3.37808
R15111 a_11023_n22908.n49 a_11023_n22908.n48 3.37783
R15112 a_11023_n22908.n43 a_11023_n22908.n1 1.89107
R15113 a_11023_n22908.n24 a_11023_n22908.n21 1.15666
R15114 a_11023_n22908.n44 a_11023_n22908.t10 0.6505
R15115 a_11023_n22908.n44 a_11023_n22908.t14 0.6505
R15116 a_11023_n22908.n46 a_11023_n22908.t13 0.6505
R15117 a_11023_n22908.n46 a_11023_n22908.t16 0.6505
R15118 a_11023_n22908.n19 a_11023_n22908.t15 0.6505
R15119 a_11023_n22908.n19 a_11023_n22908.t18 0.6505
R15120 a_11023_n22908.n18 a_11023_n22908.t17 0.6505
R15121 a_11023_n22908.n18 a_11023_n22908.t11 0.6505
R15122 a_11023_n22908.n49 a_11023_n22908.t12 0.6505
R15123 a_11023_n22908.t19 a_11023_n22908.n49 0.6505
R15124 a_11023_n22908.n38 a_11023_n22908.t7 0.5855
R15125 a_11023_n22908.n38 a_11023_n22908.t1 0.5855
R15126 a_11023_n22908.n37 a_11023_n22908.t5 0.5855
R15127 a_11023_n22908.n37 a_11023_n22908.t8 0.5855
R15128 a_11023_n22908.n36 a_11023_n22908.t2 0.5855
R15129 a_11023_n22908.n36 a_11023_n22908.t9 0.5855
R15130 a_11023_n22908.n35 a_11023_n22908.t3 0.5855
R15131 a_11023_n22908.n35 a_11023_n22908.t6 0.5855
R15132 a_11023_n22908.n34 a_11023_n22908.t0 0.5855
R15133 a_11023_n22908.n34 a_11023_n22908.t4 0.5855
R15134 a_11023_n22908.n43 a_11023_n22908.n42 0.41138
R15135 a_11023_n22908.n45 a_11023_n22908.n43 0.373278
R15136 a_11023_n22908.n40 a_11023_n22908.n39 0.183939
R15137 a_11023_n22908.n41 a_11023_n22908.n40 0.183939
R15138 a_11023_n22908.n42 a_11023_n22908.n41 0.183939
R15139 a_11023_n22908.n48 a_11023_n22908.n20 0.159616
R15140 a_11023_n22908.n48 a_11023_n22908.n47 0.159616
R15141 a_11023_n22908.n47 a_11023_n22908.n45 0.159616
R15142 a_11023_n22908.n22 a_11023_n22908.n21 0.121859
R15143 a_11023_n22908.n23 a_11023_n22908.n22 0.11975
R15144 a_11023_n22908.n17 a_11023_n22908.n2 0.11975
R15145 a_11023_n22908.n4 a_11023_n22908.n16 0.11975
R15146 a_11023_n22908.n5 a_11023_n22908.n14 0.11975
R15147 a_11023_n22908.n6 a_11023_n22908.n12 0.11975
R15148 a_11023_n22908.n25 a_11023_n22908.n24 0.11975
R15149 a_11023_n22908.n26 a_11023_n22908.n25 0.11975
R15150 a_11023_n22908.n26 a_11023_n22908.n0 0.11975
R15151 a_11023_n22908.n1 a_11023_n22908.n15 0.11975
R15152 a_11023_n22908.n32 a_11023_n22908.n15 0.11975
R15153 a_11023_n22908.n32 a_11023_n22908.n31 0.11975
R15154 a_11023_n22908.n31 a_11023_n22908.n13 0.11975
R15155 a_11023_n22908.n29 a_11023_n22908.n13 0.11975
R15156 a_11023_n22908.n29 a_11023_n22908.n28 0.11975
R15157 a_11023_n22908.n28 a_11023_n22908.n11 2.37025
R15158 a_11023_n22908.n3 a_11023_n22908.n17 0.11975
R15159 a_11023_n22908.n16 a_11023_n22908.n33 0.11975
R15160 a_11023_n22908.n14 a_11023_n22908.n30 0.11975
R15161 a_11023_n22908.n11 a_11023_n22908.n27 1.35571
R15162 a_11023_n22908.n30 a_11023_n22908.n6 0.11975
R15163 a_11023_n22908.n33 a_11023_n22908.n5 0.11975
R15164 a_11023_n22908.n4 a_11023_n22908.n3 0.11975
R15165 a_11023_n22908.n23 a_11023_n22908.n2 0.11975
R15166 a_11023_n22908.n1 a_11023_n22908.n0 0.11975
R15167 a_11023_n22908.n9 a_11023_n22908.n10 0.0946176
R15168 a_11023_n22908.n7 a_11023_n22908.n9 0.0946176
R15169 a_11023_n22908.n8 a_11023_n22908.n7 0.0946176
R15170 a_11023_n22908.n27 a_11023_n22908.n8 0.0946176
R15171 a_38256_1564.n10 a_38256_1564.t8 15.8415
R15172 a_38256_1564.n4 a_38256_1564.t17 15.8415
R15173 a_38256_1564.n5 a_38256_1564.t20 15.8415
R15174 a_38256_1564.n6 a_38256_1564.t23 15.8415
R15175 a_38256_1564.n7 a_38256_1564.t11 15.8415
R15176 a_38256_1564.n8 a_38256_1564.t14 15.8415
R15177 a_38256_1564.n9 a_38256_1564.t18 15.8415
R15178 a_38256_1564.n11 a_38256_1564.t22 15.8415
R15179 a_38256_1564.n10 a_38256_1564.t21 13.4447
R15180 a_38256_1564.n4 a_38256_1564.t12 13.4447
R15181 a_38256_1564.n5 a_38256_1564.t15 13.4447
R15182 a_38256_1564.n6 a_38256_1564.t19 13.4447
R15183 a_38256_1564.n7 a_38256_1564.t9 13.4447
R15184 a_38256_1564.n8 a_38256_1564.t10 13.4447
R15185 a_38256_1564.n9 a_38256_1564.t13 13.4447
R15186 a_38256_1564.n11 a_38256_1564.t16 13.4447
R15187 a_38256_1564.n5 a_38256_1564.n4 10.5449
R15188 a_38256_1564.n6 a_38256_1564.n5 10.5449
R15189 a_38256_1564.n7 a_38256_1564.n6 10.5449
R15190 a_38256_1564.n8 a_38256_1564.n7 10.5449
R15191 a_38256_1564.n9 a_38256_1564.n8 10.5449
R15192 a_38256_1564.n11 a_38256_1564.n9 10.5449
R15193 a_38256_1564.n11 a_38256_1564.n10 10.5449
R15194 a_38256_1564.n0 a_38256_1564.n3 7.22489
R15195 a_38256_1564.n0 a_38256_1564.n2 6.36702
R15196 a_38256_1564.n12 a_38256_1564.n0 3.56115
R15197 a_38256_1564.n0 a_38256_1564.n1 2.68463
R15198 a_38256_1564.n0 a_38256_1564.n11 2.37315
R15199 a_38256_1564.n1 a_38256_1564.t6 2.06607
R15200 a_38256_1564.t7 a_38256_1564.n12 2.06607
R15201 a_38256_1564.n3 a_38256_1564.t0 1.99806
R15202 a_38256_1564.n3 a_38256_1564.t1 1.99806
R15203 a_38256_1564.n2 a_38256_1564.t3 1.99806
R15204 a_38256_1564.n2 a_38256_1564.t2 1.99806
R15205 a_38256_1564.n1 a_38256_1564.t5 1.4923
R15206 a_38256_1564.n12 a_38256_1564.t4 1.4923
R15207 a_26553_377.n2 a_26553_377.n0 38.9364
R15208 a_26553_377.n1 a_26553_377.t5 29.2005
R15209 a_26553_377.n0 a_26553_377.t2 20.1607
R15210 a_26553_377.n2 a_26553_377.n1 17.6316
R15211 a_26553_377.n1 a_26553_377.t3 12.1428
R15212 a_26553_377.n3 a_26553_377.n2 11.8939
R15213 a_26553_377.n0 a_26553_377.t4 10.8288
R15214 a_26553_377.n3 a_26553_377.t0 8.67092
R15215 a_26553_377.t1 a_26553_377.n3 4.67457
R15216 a_33496_n6659.n6 a_33496_n6659.t28 15.4765
R15217 a_33496_n6659.n7 a_33496_n6659.t25 15.4765
R15218 a_33496_n6659.n8 a_33496_n6659.t30 15.4765
R15219 a_33496_n6659.n9 a_33496_n6659.t32 15.4765
R15220 a_33496_n6659.n10 a_33496_n6659.t39 15.4765
R15221 a_33496_n6659.n11 a_33496_n6659.t12 15.4765
R15222 a_33496_n6659.n12 a_33496_n6659.t8 15.4765
R15223 a_33496_n6659.n13 a_33496_n6659.t9 15.4765
R15224 a_33496_n6659.n14 a_33496_n6659.t22 15.4765
R15225 a_33496_n6659.n15 a_33496_n6659.t18 15.4765
R15226 a_33496_n6659.n1 a_33496_n6659.t24 15.4765
R15227 a_33496_n6659.n2 a_33496_n6659.t19 15.4765
R15228 a_33496_n6659.n3 a_33496_n6659.t38 15.4765
R15229 a_33496_n6659.n4 a_33496_n6659.t34 15.4765
R15230 a_33496_n6659.n5 a_33496_n6659.t37 15.4765
R15231 a_33496_n6659.n0 a_33496_n6659.t33 15.4765
R15232 a_33496_n6659.n0 a_33496_n6659.t3 14.6183
R15233 a_33496_n6659.n6 a_33496_n6659.t10 11.863
R15234 a_33496_n6659.n7 a_33496_n6659.t16 11.863
R15235 a_33496_n6659.n8 a_33496_n6659.t20 11.863
R15236 a_33496_n6659.n9 a_33496_n6659.t21 11.863
R15237 a_33496_n6659.n10 a_33496_n6659.t17 11.863
R15238 a_33496_n6659.n11 a_33496_n6659.t35 11.863
R15239 a_33496_n6659.n12 a_33496_n6659.t29 11.863
R15240 a_33496_n6659.n13 a_33496_n6659.t31 11.863
R15241 a_33496_n6659.n14 a_33496_n6659.t36 11.863
R15242 a_33496_n6659.n15 a_33496_n6659.t11 11.863
R15243 a_33496_n6659.n3 a_33496_n6659.t27 11.863
R15244 a_33496_n6659.n4 a_33496_n6659.t23 11.863
R15245 a_33496_n6659.n5 a_33496_n6659.t26 11.863
R15246 a_33496_n6659.n0 a_33496_n6659.t14 11.863
R15247 a_33496_n6659.n1 a_33496_n6659.t15 11.8022
R15248 a_33496_n6659.n2 a_33496_n6659.t13 11.8022
R15249 a_33496_n6659.n0 a_33496_n6659.t1 11.3584
R15250 a_33496_n6659.n7 a_33496_n6659.n6 10.5449
R15251 a_33496_n6659.n8 a_33496_n6659.n7 10.5449
R15252 a_33496_n6659.n9 a_33496_n6659.n8 10.5449
R15253 a_33496_n6659.n10 a_33496_n6659.n9 10.5449
R15254 a_33496_n6659.n11 a_33496_n6659.n10 10.5449
R15255 a_33496_n6659.n12 a_33496_n6659.n11 10.5449
R15256 a_33496_n6659.n13 a_33496_n6659.n12 10.5449
R15257 a_33496_n6659.n14 a_33496_n6659.n13 10.5449
R15258 a_33496_n6659.n15 a_33496_n6659.n14 10.5449
R15259 a_33496_n6659.n1 a_33496_n6659.n15 10.5449
R15260 a_33496_n6659.n4 a_33496_n6659.n3 10.5449
R15261 a_33496_n6659.n5 a_33496_n6659.n4 10.5449
R15262 a_33496_n6659.n0 a_33496_n6659.n5 10.5449
R15263 a_33496_n6659.n0 a_33496_n6659.n2 10.5449
R15264 a_33496_n6659.n0 a_33496_n6659.t7 10.4819
R15265 a_33496_n6659.n0 a_33496_n6659.t0 10.4819
R15266 a_33496_n6659.n0 a_33496_n6659.t6 10.4819
R15267 a_33496_n6659.n2 a_33496_n6659.n1 10.3816
R15268 a_33496_n6659.n0 a_33496_n6659.t5 9.32628
R15269 a_33496_n6659.n0 a_33496_n6659.t4 8.44976
R15270 a_33496_n6659.t2 a_33496_n6659.n0 8.44976
R15271 a_31628_n5940.n26 a_31628_n5940.t39 31.6987
R15272 a_31628_n5940.n24 a_31628_n5940.t36 31.6987
R15273 a_31628_n5940.n27 a_31628_n5940.t41 18.6885
R15274 a_31628_n5940.n28 a_31628_n5940.t37 18.6885
R15275 a_31628_n5940.n26 a_31628_n5940.t45 18.6885
R15276 a_31628_n5940.n24 a_31628_n5940.t42 18.6885
R15277 a_31628_n5940.n22 a_31628_n5940.t32 18.6885
R15278 a_31628_n5940.n23 a_31628_n5940.t35 18.6885
R15279 a_31628_n5940.n30 a_31628_n5940.n25 17.1811
R15280 a_31628_n5940.n27 a_31628_n5940.t40 11.133
R15281 a_31628_n5940.n28 a_31628_n5940.t43 11.133
R15282 a_31628_n5940.n26 a_31628_n5940.t44 11.133
R15283 a_31628_n5940.n24 a_31628_n5940.t33 11.133
R15284 a_31628_n5940.n22 a_31628_n5940.t38 11.133
R15285 a_31628_n5940.n23 a_31628_n5940.t34 11.133
R15286 a_31628_n5940.n28 a_31628_n5940.n27 10.5449
R15287 a_31628_n5940.n23 a_31628_n5940.n22 10.5449
R15288 a_31628_n5940.n19 a_31628_n5940.n18 7.0655
R15289 a_31628_n5940.n13 a_31628_n5940.n12 7.0655
R15290 a_31628_n5940.n29 a_31628_n5940.n26 6.48939
R15291 a_31628_n5940.n25 a_31628_n5940.n24 6.48939
R15292 a_31628_n5940.n2 a_31628_n5940.n15 6.4355
R15293 a_31628_n5940.n20 a_31628_n5940.n16 6.4355
R15294 a_31628_n5940.n19 a_31628_n5940.n17 6.4355
R15295 a_31628_n5940.n13 a_31628_n5940.n11 6.4355
R15296 a_31628_n5940.n14 a_31628_n5940.n10 6.4355
R15297 a_31628_n5940.n1 a_31628_n5940.n9 6.4355
R15298 a_31628_n5940.n30 a_31628_n5940.n29 6.02113
R15299 a_31628_n5940.n31 a_31628_n5940.n30 5.5805
R15300 a_31628_n5940.n29 a_31628_n5940.n28 4.05606
R15301 a_31628_n5940.n25 a_31628_n5940.n23 4.05606
R15302 a_31628_n5940.n15 a_31628_n5940.t14 3.37782
R15303 a_31628_n5940.n15 a_31628_n5940.t0 3.37782
R15304 a_31628_n5940.n16 a_31628_n5940.t13 3.37782
R15305 a_31628_n5940.n16 a_31628_n5940.t11 3.37782
R15306 a_31628_n5940.n17 a_31628_n5940.t5 3.37782
R15307 a_31628_n5940.n17 a_31628_n5940.t12 3.37782
R15308 a_31628_n5940.n18 a_31628_n5940.t4 3.37782
R15309 a_31628_n5940.n18 a_31628_n5940.t6 3.37782
R15310 a_31628_n5940.n12 a_31628_n5940.t10 3.37782
R15311 a_31628_n5940.n12 a_31628_n5940.t15 3.37782
R15312 a_31628_n5940.n11 a_31628_n5940.t7 3.37782
R15313 a_31628_n5940.n11 a_31628_n5940.t8 3.37782
R15314 a_31628_n5940.n10 a_31628_n5940.t1 3.37782
R15315 a_31628_n5940.n10 a_31628_n5940.t9 3.37782
R15316 a_31628_n5940.n9 a_31628_n5940.t2 3.37782
R15317 a_31628_n5940.n9 a_31628_n5940.t3 3.37782
R15318 a_31628_n5940.n5 a_31628_n5940.n3 2.93257
R15319 a_31628_n5940.n31 a_31628_n5940.n21 2.62533
R15320 a_31628_n5940.n5 a_31628_n5940.n4 2.6005
R15321 a_31628_n5940.n7 a_31628_n5940.n6 2.6005
R15322 a_31628_n5940.n0 a_31628_n5940.n8 2.6005
R15323 a_31628_n5940.n35 a_31628_n5940.n34 2.6005
R15324 a_31628_n5940.n33 a_31628_n5940.n32 2.6005
R15325 a_31628_n5940.n36 a_31628_n5940.n1 2.6005
R15326 a_31628_n5940.n21 a_31628_n5940.t23 2.06607
R15327 a_31628_n5940.n32 a_31628_n5940.t22 2.06607
R15328 a_31628_n5940.n34 a_31628_n5940.t16 2.06607
R15329 a_31628_n5940.n8 a_31628_n5940.t26 2.06607
R15330 a_31628_n5940.n6 a_31628_n5940.t25 2.06607
R15331 a_31628_n5940.n4 a_31628_n5940.t20 2.06607
R15332 a_31628_n5940.n3 a_31628_n5940.t17 2.06607
R15333 a_31628_n5940.t31 a_31628_n5940.n36 2.06607
R15334 a_31628_n5940.n21 a_31628_n5940.t24 1.4923
R15335 a_31628_n5940.n32 a_31628_n5940.t21 1.4923
R15336 a_31628_n5940.n34 a_31628_n5940.t29 1.4923
R15337 a_31628_n5940.n8 a_31628_n5940.t28 1.4923
R15338 a_31628_n5940.n6 a_31628_n5940.t27 1.4923
R15339 a_31628_n5940.n4 a_31628_n5940.t18 1.4923
R15340 a_31628_n5940.n3 a_31628_n5940.t19 1.4923
R15341 a_31628_n5940.n36 a_31628_n5940.t30 1.4923
R15342 a_31628_n5940.n1 a_31628_n5940.n14 0.6305
R15343 a_31628_n5940.n14 a_31628_n5940.n13 0.6305
R15344 a_31628_n5940.n20 a_31628_n5940.n19 0.6305
R15345 a_31628_n5940.n2 a_31628_n5940.n20 0.6305
R15346 a_31628_n5940.n1 a_31628_n5940.n0 0.4039
R15347 a_31628_n5940.n7 a_31628_n5940.n5 0.348086
R15348 a_31628_n5940.n0 a_31628_n5940.n7 0.348086
R15349 a_31628_n5940.n1 a_31628_n5940.n35 0.348086
R15350 a_31628_n5940.n35 a_31628_n5940.n33 0.348086
R15351 a_31628_n5940.n33 a_31628_n5940.n31 0.323259
R15352 a_31628_n5940.n1 a_31628_n5940.n2 0.315406
R15353 a_27884_332.n2 a_27884_332.n0 37.0046
R15354 a_27884_332.n1 a_27884_332.t2 21.499
R15355 a_27884_332.n2 a_27884_332.n1 20.7028
R15356 a_27884_332.n0 a_27884_332.t3 18.9805
R15357 a_27884_332.t1 a_27884_332.n2 13.073
R15358 a_27884_332.n0 a_27884_332.t5 11.4372
R15359 a_27884_332.t1 a_27884_332.t0 8.92356
R15360 a_27884_332.n1 a_27884_332.t4 8.69967
R15361 a_29800_n5940.n5 a_29800_n5940.t19 15.7685
R15362 a_29800_n5940.n6 a_29800_n5940.t17 15.7685
R15363 a_29800_n5940.n7 a_29800_n5940.t10 15.7685
R15364 a_29800_n5940.n8 a_29800_n5940.t18 15.7685
R15365 a_29800_n5940.n9 a_29800_n5940.t11 15.7685
R15366 a_29800_n5940.n10 a_29800_n5940.t8 15.7685
R15367 a_29800_n5940.n3 a_29800_n5940.t9 15.7685
R15368 a_29800_n5940.n4 a_29800_n5940.t14 15.7685
R15369 a_29800_n5940.n5 a_29800_n5940.t7 11.6197
R15370 a_29800_n5940.n6 a_29800_n5940.t12 11.6197
R15371 a_29800_n5940.n7 a_29800_n5940.t15 11.6197
R15372 a_29800_n5940.n8 a_29800_n5940.t13 11.6197
R15373 a_29800_n5940.n9 a_29800_n5940.t16 11.6197
R15374 a_29800_n5940.n10 a_29800_n5940.t20 11.6197
R15375 a_29800_n5940.n3 a_29800_n5940.t22 11.6197
R15376 a_29800_n5940.n4 a_29800_n5940.t21 11.6197
R15377 a_29800_n5940.n6 a_29800_n5940.n5 10.5449
R15378 a_29800_n5940.n7 a_29800_n5940.n6 10.5449
R15379 a_29800_n5940.n8 a_29800_n5940.n7 10.5449
R15380 a_29800_n5940.n9 a_29800_n5940.n8 10.5449
R15381 a_29800_n5940.n10 a_29800_n5940.n9 10.5449
R15382 a_29800_n5940.n4 a_29800_n5940.n3 10.5449
R15383 a_29800_n5940.n0 a_29800_n5940.t2 10.4819
R15384 a_29800_n5940.n11 a_29800_n5940.n10 8.41578
R15385 a_29800_n5940.n0 a_29800_n5940.n2 7.31398
R15386 a_29800_n5940.n12 a_29800_n5940.n0 6.25311
R15387 a_29800_n5940.n0 a_29800_n5940.n1 5.37659
R15388 a_29800_n5940.n2 a_29800_n5940.t0 4.04494
R15389 a_29800_n5940.n2 a_29800_n5940.t1 4.04494
R15390 a_29800_n5940.n1 a_29800_n5940.t3 3.07367
R15391 a_29800_n5940.n1 a_29800_n5940.t4 3.07367
R15392 a_29800_n5940.t6 a_29800_n5940.n12 3.07367
R15393 a_29800_n5940.n12 a_29800_n5940.t5 3.07367
R15394 a_29800_n5940.n0 a_29800_n5940.n11 2.93567
R15395 a_29800_n5940.n11 a_29800_n5940.n4 2.12967
R15396 a_28156_n6412.n8 a_28156_n6412.t21 31.6987
R15397 a_28156_n6412.n12 a_28156_n6412.t23 31.6987
R15398 a_28156_n6412.n8 a_28156_n6412.t17 18.6885
R15399 a_28156_n6412.n6 a_28156_n6412.t18 18.6885
R15400 a_28156_n6412.n7 a_28156_n6412.t27 18.6885
R15401 a_28156_n6412.n12 a_28156_n6412.t19 18.6885
R15402 a_28156_n6412.n10 a_28156_n6412.t24 18.6885
R15403 a_28156_n6412.n11 a_28156_n6412.t28 18.6885
R15404 a_28156_n6412.n0 a_28156_n6412.n14 15.1205
R15405 a_28156_n6412.n12 a_28156_n6412.t22 11.1938
R15406 a_28156_n6412.n10 a_28156_n6412.t16 11.1938
R15407 a_28156_n6412.n11 a_28156_n6412.t29 11.1938
R15408 a_28156_n6412.n8 a_28156_n6412.t20 11.133
R15409 a_28156_n6412.n6 a_28156_n6412.t25 11.133
R15410 a_28156_n6412.n7 a_28156_n6412.t26 11.133
R15411 a_28156_n6412.n7 a_28156_n6412.n6 10.5449
R15412 a_28156_n6412.n11 a_28156_n6412.n10 10.5449
R15413 a_28156_n6412.n14 a_28156_n6412.n13 7.23613
R15414 a_28156_n6412.n2 a_28156_n6412.n18 7.13263
R15415 a_28156_n6412.n1 a_28156_n6412.n16 7.13263
R15416 a_28156_n6412.n9 a_28156_n6412.n8 6.48939
R15417 a_28156_n6412.n13 a_28156_n6412.n12 6.48939
R15418 a_28156_n6412.n2 a_28156_n6412.n17 6.43746
R15419 a_28156_n6412.n1 a_28156_n6412.n15 6.43746
R15420 a_28156_n6412.n14 a_28156_n6412.n9 6.15613
R15421 a_28156_n6412.n9 a_28156_n6412.n7 4.05606
R15422 a_28156_n6412.n13 a_28156_n6412.n11 4.05606
R15423 a_28156_n6412.n18 a_28156_n6412.t0 3.8098
R15424 a_28156_n6412.n18 a_28156_n6412.t1 3.8098
R15425 a_28156_n6412.n17 a_28156_n6412.t2 3.8098
R15426 a_28156_n6412.n17 a_28156_n6412.t3 3.8098
R15427 a_28156_n6412.n15 a_28156_n6412.t5 3.8098
R15428 a_28156_n6412.n15 a_28156_n6412.t4 3.8098
R15429 a_28156_n6412.n16 a_28156_n6412.t6 3.8098
R15430 a_28156_n6412.n16 a_28156_n6412.t7 3.8098
R15431 a_28156_n6412.n0 a_28156_n6412.n3 3.34593
R15432 a_28156_n6412.n0 a_28156_n6412.n5 2.78906
R15433 a_28156_n6412.n0 a_28156_n6412.n4 2.71593
R15434 a_28156_n6412.n19 a_28156_n6412.n0 2.71593
R15435 a_28156_n6412.n5 a_28156_n6412.t10 2.06607
R15436 a_28156_n6412.n5 a_28156_n6412.t8 2.06607
R15437 a_28156_n6412.n4 a_28156_n6412.t9 2.06607
R15438 a_28156_n6412.n4 a_28156_n6412.t13 2.06607
R15439 a_28156_n6412.n3 a_28156_n6412.t14 2.06607
R15440 a_28156_n6412.n3 a_28156_n6412.t11 2.06607
R15441 a_28156_n6412.t15 a_28156_n6412.n19 2.06607
R15442 a_28156_n6412.n19 a_28156_n6412.t12 2.06607
R15443 a_28156_n6412.n0 a_28156_n6412.n1 1.35405
R15444 a_28156_n6412.n1 a_28156_n6412.n2 0.577741
R15445 a_11023_n12196.n2 a_11023_n12196.t38 56.019
R15446 a_11023_n12196.n1 a_11023_n12196.t26 55.9719
R15447 a_11023_n12196.n1 a_11023_n12196.t34 55.9719
R15448 a_11023_n12196.n1 a_11023_n12196.t21 55.9719
R15449 a_11023_n12196.n1 a_11023_n12196.t36 55.9719
R15450 a_11023_n12196.n1 a_11023_n12196.t23 55.9719
R15451 a_11023_n12196.n1 a_11023_n12196.t30 55.9719
R15452 a_11023_n12196.n1 a_11023_n12196.t39 55.9719
R15453 a_11023_n12196.n1 a_11023_n12196.t25 55.9719
R15454 a_11023_n12196.n1 a_11023_n12196.t31 55.9719
R15455 a_11023_n12196.n2 a_11023_n12196.t27 55.9719
R15456 a_11023_n12196.n2 a_11023_n12196.t33 55.9719
R15457 a_11023_n12196.n2 a_11023_n12196.t20 55.9719
R15458 a_11023_n12196.n2 a_11023_n12196.t28 55.9719
R15459 a_11023_n12196.n2 a_11023_n12196.t35 55.9719
R15460 a_11023_n12196.n2 a_11023_n12196.t22 55.9719
R15461 a_11023_n12196.n2 a_11023_n12196.t37 55.9719
R15462 a_11023_n12196.n2 a_11023_n12196.t24 55.9719
R15463 a_11023_n12196.n2 a_11023_n12196.t32 55.9719
R15464 a_11023_n12196.n1 a_11023_n12196.n0 0.14323
R15465 a_11023_n12196.n3 a_11023_n12196.t16 3.87048
R15466 a_11023_n12196.n3 a_11023_n12196.t0 3.68704
R15467 a_11023_n12196.n4 a_11023_n12196.t6 3.68704
R15468 a_11023_n12196.n5 a_11023_n12196.t2 3.68704
R15469 a_11023_n12196.n6 a_11023_n12196.t8 3.68704
R15470 a_11023_n12196.n11 a_11023_n12196.t18 3.53719
R15471 a_11023_n12196.n8 a_11023_n12196.t11 3.37808
R15472 a_11023_n12196.n9 a_11023_n12196.t5 3.37808
R15473 a_11023_n12196.n10 a_11023_n12196.t9 3.37808
R15474 a_11023_n12196.t15 a_11023_n12196.n11 3.37783
R15475 a_11023_n12196.t11 a_11023_n12196.t4 0.6505
R15476 a_11023_n12196.t5 a_11023_n12196.t19 0.6505
R15477 a_11023_n12196.t9 a_11023_n12196.t14 0.6505
R15478 a_11023_n12196.t18 a_11023_n12196.t10 0.6505
R15479 a_11023_n12196.t3 a_11023_n12196.t15 0.6505
R15480 a_11023_n12196.t16 a_11023_n12196.t7 0.5855
R15481 a_11023_n12196.t0 a_11023_n12196.t13 0.5855
R15482 a_11023_n12196.t6 a_11023_n12196.t12 0.5855
R15483 a_11023_n12196.t2 a_11023_n12196.t17 0.5855
R15484 a_11023_n12196.t8 a_11023_n12196.t1 0.5855
R15485 a_11023_n12196.n7 a_11023_n12196.n6 0.41138
R15486 a_11023_n12196.n8 a_11023_n12196.n7 0.373278
R15487 a_11023_n12196.n4 a_11023_n12196.n3 0.183939
R15488 a_11023_n12196.n5 a_11023_n12196.n4 0.183939
R15489 a_11023_n12196.n6 a_11023_n12196.n5 0.183939
R15490 a_11023_n12196.n11 a_11023_n12196.n10 0.159616
R15491 a_11023_n12196.n10 a_11023_n12196.n9 0.159616
R15492 a_11023_n12196.n9 a_11023_n12196.n8 0.159616
R15493 a_11023_n12196.n1 a_11023_n12196.t29 56.3117
R15494 a_11023_n12196.n7 a_11023_n12196.n0 2.08751
R15495 a_11023_n12196.n0 a_11023_n12196.n2 2.43655
R15496 a_11087_n12816.n26 a_11087_n12816.t30 14.9789
R15497 a_11087_n12816.n11 a_11087_n12816.n9 10.553
R15498 a_11087_n12816.n26 a_11087_n12816.n25 10.4369
R15499 a_11087_n12816.n28 a_11087_n12816.n27 10.4369
R15500 a_11087_n12816.n24 a_11087_n12816.n23 10.4308
R15501 a_11087_n12816.n22 a_11087_n12816.n21 10.4308
R15502 a_11087_n12816.n20 a_11087_n12816.n19 10.4308
R15503 a_11087_n12816.n11 a_11087_n12816.n10 10.4156
R15504 a_11087_n12816.n15 a_11087_n12816.n14 10.4129
R15505 a_11087_n12816.n17 a_11087_n12816.n16 10.4121
R15506 a_11087_n12816.n13 a_11087_n12816.n12 10.4121
R15507 a_11087_n12816.n2 a_11087_n12816.n0 10.357
R15508 a_11087_n12816.n8 a_11087_n12816.n7 10.2004
R15509 a_11087_n12816.n4 a_11087_n12816.n3 10.2004
R15510 a_11087_n12816.n6 a_11087_n12816.n5 10.198
R15511 a_11087_n12816.n2 a_11087_n12816.n1 10.1921
R15512 a_11087_n12816.n18 a_11087_n12816.n8 0.773592
R15513 a_11087_n12816.n7 a_11087_n12816.t12 0.6505
R15514 a_11087_n12816.n7 a_11087_n12816.t16 0.6505
R15515 a_11087_n12816.n5 a_11087_n12816.t11 0.6505
R15516 a_11087_n12816.n5 a_11087_n12816.t19 0.6505
R15517 a_11087_n12816.n3 a_11087_n12816.t14 0.6505
R15518 a_11087_n12816.n3 a_11087_n12816.t18 0.6505
R15519 a_11087_n12816.n1 a_11087_n12816.t17 0.6505
R15520 a_11087_n12816.n1 a_11087_n12816.t10 0.6505
R15521 a_11087_n12816.n0 a_11087_n12816.t15 0.6505
R15522 a_11087_n12816.n0 a_11087_n12816.t13 0.6505
R15523 a_11087_n12816.n25 a_11087_n12816.t6 0.5855
R15524 a_11087_n12816.n25 a_11087_n12816.t0 0.5855
R15525 a_11087_n12816.n23 a_11087_n12816.t2 0.5855
R15526 a_11087_n12816.n23 a_11087_n12816.t5 0.5855
R15527 a_11087_n12816.n21 a_11087_n12816.t1 0.5855
R15528 a_11087_n12816.n21 a_11087_n12816.t8 0.5855
R15529 a_11087_n12816.n19 a_11087_n12816.t4 0.5855
R15530 a_11087_n12816.n19 a_11087_n12816.t7 0.5855
R15531 a_11087_n12816.n16 a_11087_n12816.t26 0.5855
R15532 a_11087_n12816.n16 a_11087_n12816.t22 0.5855
R15533 a_11087_n12816.n14 a_11087_n12816.t27 0.5855
R15534 a_11087_n12816.n14 a_11087_n12816.t29 0.5855
R15535 a_11087_n12816.n12 a_11087_n12816.t24 0.5855
R15536 a_11087_n12816.n12 a_11087_n12816.t20 0.5855
R15537 a_11087_n12816.n10 a_11087_n12816.t21 0.5855
R15538 a_11087_n12816.n10 a_11087_n12816.t28 0.5855
R15539 a_11087_n12816.n9 a_11087_n12816.t23 0.5855
R15540 a_11087_n12816.n9 a_11087_n12816.t25 0.5855
R15541 a_11087_n12816.t9 a_11087_n12816.n28 0.5855
R15542 a_11087_n12816.n28 a_11087_n12816.t3 0.5855
R15543 a_11087_n12816.n18 a_11087_n12816.n17 0.366893
R15544 a_11087_n12816.n20 a_11087_n12816.n18 0.297718
R15545 a_11087_n12816.n27 a_11087_n12816.n26 0.1615
R15546 a_11087_n12816.n8 a_11087_n12816.n6 0.161
R15547 a_11087_n12816.n4 a_11087_n12816.n2 0.1605
R15548 a_11087_n12816.n6 a_11087_n12816.n4 0.1605
R15549 a_11087_n12816.n22 a_11087_n12816.n20 0.1605
R15550 a_11087_n12816.n24 a_11087_n12816.n22 0.1605
R15551 a_11087_n12816.n27 a_11087_n12816.n24 0.1585
R15552 a_11087_n12816.n17 a_11087_n12816.n15 0.139126
R15553 a_11087_n12816.n13 a_11087_n12816.n11 0.136566
R15554 a_11087_n12816.n15 a_11087_n12816.n13 0.13486
R15555 a_21772_n20836.n5 a_21772_n20836.t20 15.8415
R15556 a_21772_n20836.n6 a_21772_n20836.t23 15.8415
R15557 a_21772_n20836.n7 a_21772_n20836.t9 15.8415
R15558 a_21772_n20836.n8 a_21772_n20836.t21 15.8415
R15559 a_21772_n20836.n9 a_21772_n20836.t18 15.8415
R15560 a_21772_n20836.n10 a_21772_n20836.t19 15.8415
R15561 a_21772_n20836.n4 a_21772_n20836.t8 15.8415
R15562 a_21772_n20836.n11 a_21772_n20836.t22 15.8415
R15563 a_21772_n20836.n5 a_21772_n20836.t13 13.4447
R15564 a_21772_n20836.n6 a_21772_n20836.t10 13.4447
R15565 a_21772_n20836.n7 a_21772_n20836.t17 13.4447
R15566 a_21772_n20836.n8 a_21772_n20836.t14 13.4447
R15567 a_21772_n20836.n9 a_21772_n20836.t11 13.4447
R15568 a_21772_n20836.n10 a_21772_n20836.t12 13.4447
R15569 a_21772_n20836.n4 a_21772_n20836.t16 13.4447
R15570 a_21772_n20836.n11 a_21772_n20836.t15 13.4447
R15571 a_21772_n20836.n6 a_21772_n20836.n5 10.5449
R15572 a_21772_n20836.n7 a_21772_n20836.n6 10.5449
R15573 a_21772_n20836.n8 a_21772_n20836.n7 10.5449
R15574 a_21772_n20836.n9 a_21772_n20836.n8 10.5449
R15575 a_21772_n20836.n10 a_21772_n20836.n9 10.5449
R15576 a_21772_n20836.n11 a_21772_n20836.n4 10.5449
R15577 a_21772_n20836.n11 a_21772_n20836.n10 10.5449
R15578 a_21772_n20836.n0 a_21772_n20836.n3 7.22489
R15579 a_21772_n20836.n0 a_21772_n20836.n2 6.36702
R15580 a_21772_n20836.n12 a_21772_n20836.n0 3.56115
R15581 a_21772_n20836.n0 a_21772_n20836.n1 2.68463
R15582 a_21772_n20836.n0 a_21772_n20836.n11 2.37183
R15583 a_21772_n20836.n1 a_21772_n20836.t5 2.06607
R15584 a_21772_n20836.t7 a_21772_n20836.n12 2.06607
R15585 a_21772_n20836.n2 a_21772_n20836.t3 1.99806
R15586 a_21772_n20836.n2 a_21772_n20836.t2 1.99806
R15587 a_21772_n20836.n3 a_21772_n20836.t1 1.99806
R15588 a_21772_n20836.n3 a_21772_n20836.t0 1.99806
R15589 a_21772_n20836.n1 a_21772_n20836.t6 1.4923
R15590 a_21772_n20836.n12 a_21772_n20836.t4 1.4923
R15591 a_13623_n6840.n1 a_13623_n6840.t30 56.1018
R15592 a_13623_n6840.n2 a_13623_n6840.t39 56.0719
R15593 a_13623_n6840.n1 a_13623_n6840.t17 56.0141
R15594 a_13623_n6840.n1 a_13623_n6840.t25 55.9719
R15595 a_13623_n6840.n1 a_13623_n6840.t37 55.9719
R15596 a_13623_n6840.n1 a_13623_n6840.t32 55.9719
R15597 a_13623_n6840.n1 a_13623_n6840.t44 55.9719
R15598 a_13623_n6840.n1 a_13623_n6840.t34 55.9719
R15599 a_13623_n6840.n1 a_13623_n6840.t29 55.9719
R15600 a_13623_n6840.n1 a_13623_n6840.t41 55.9719
R15601 a_13623_n6840.n1 a_13623_n6840.t36 55.9719
R15602 a_13623_n6840.n1 a_13623_n6840.t20 55.9719
R15603 a_13623_n6840.n1 a_13623_n6840.t40 55.9719
R15604 a_13623_n6840.n1 a_13623_n6840.t27 55.9719
R15605 a_13623_n6840.n1 a_13623_n6840.t19 55.9719
R15606 a_13623_n6840.n1 a_13623_n6840.t33 55.9719
R15607 a_13623_n6840.n1 a_13623_n6840.t23 55.9719
R15608 a_13623_n6840.n1 a_13623_n6840.t16 55.9719
R15609 a_13623_n6840.n1 a_13623_n6840.t31 55.9719
R15610 a_13623_n6840.n1 a_13623_n6840.t26 55.9719
R15611 a_13623_n6840.n1 a_13623_n6840.t38 55.9719
R15612 a_13623_n6840.n2 a_13623_n6840.t22 55.9719
R15613 a_13623_n6840.n2 a_13623_n6840.t45 55.9719
R15614 a_13623_n6840.n2 a_13623_n6840.t35 55.9719
R15615 a_13623_n6840.n2 a_13623_n6840.t18 55.9719
R15616 a_13623_n6840.n2 a_13623_n6840.t42 55.9719
R15617 a_13623_n6840.n2 a_13623_n6840.t28 55.9719
R15618 a_13623_n6840.n4 a_13623_n6840.t21 55.9719
R15619 a_13623_n6840.n4 a_13623_n6840.t43 55.9719
R15620 a_13623_n6840.n4 a_13623_n6840.t24 55.9719
R15621 a_13623_n6840.n0 a_13623_n6840.n1 46.1399
R15622 a_13623_n6840.n0 a_13623_n6840.n9 6.90733
R15623 a_13623_n6840.n3 a_13623_n6840.n11 6.89497
R15624 a_13623_n6840.n3 a_13623_n6840.n10 6.3768
R15625 a_13623_n6840.n0 a_13623_n6840.n8 6.3768
R15626 a_13623_n6840.n12 a_13623_n6840.n0 3.21104
R15627 a_13623_n6840.n0 a_13623_n6840.n6 2.7042
R15628 a_13623_n6840.n0 a_13623_n6840.n7 2.7042
R15629 a_13623_n6840.n0 a_13623_n6840.n5 2.7042
R15630 a_13623_n6840.n6 a_13623_n6840.t14 2.06607
R15631 a_13623_n6840.n7 a_13623_n6840.t11 2.06607
R15632 a_13623_n6840.n5 a_13623_n6840.t13 2.06607
R15633 a_13623_n6840.t15 a_13623_n6840.n12 2.06607
R15634 a_13623_n6840.n10 a_13623_n6840.t5 1.99806
R15635 a_13623_n6840.n10 a_13623_n6840.t6 1.99806
R15636 a_13623_n6840.n11 a_13623_n6840.t1 1.99806
R15637 a_13623_n6840.n11 a_13623_n6840.t2 1.99806
R15638 a_13623_n6840.n9 a_13623_n6840.t7 1.99806
R15639 a_13623_n6840.n9 a_13623_n6840.t4 1.99806
R15640 a_13623_n6840.n8 a_13623_n6840.t3 1.99806
R15641 a_13623_n6840.n8 a_13623_n6840.t0 1.99806
R15642 a_13623_n6840.n6 a_13623_n6840.t10 1.4923
R15643 a_13623_n6840.n7 a_13623_n6840.t8 1.4923
R15644 a_13623_n6840.n5 a_13623_n6840.t12 1.4923
R15645 a_13623_n6840.n12 a_13623_n6840.t9 1.4923
R15646 a_13623_n6840.n0 a_13623_n6840.n3 1.35826
R15647 a_13623_n6840.n1 a_13623_n6840.n4 1.21355
R15648 a_13623_n6840.n4 a_13623_n6840.n2 0.8005
R15649 a_21692_n6694.n8 a_21692_n6694.n6 23.6386
R15650 a_21692_n6694.n1 a_21692_n6694.n24 23.1113
R15651 a_21692_n6694.n12 a_21692_n6694.t5 20.0755
R15652 a_21692_n6694.n27 a_21692_n6694.t30 19.5645
R15653 a_21692_n6694.n25 a_21692_n6694.t4 18.6885
R15654 a_21692_n6694.n3 a_21692_n6694.t34 18.6885
R15655 a_21692_n6694.n12 a_21692_n6694.t31 18.3519
R15656 a_21692_n6694.n8 a_21692_n6694.n7 17.9041
R15657 a_21692_n6694.n18 a_21692_n6694.t7 17.7395
R15658 a_21692_n6694.n13 a_21692_n6694.t27 17.3502
R15659 a_21692_n6694.n27 a_21692_n6694.t22 17.1312
R15660 a_21692_n6694.n30 a_21692_n6694.n4 17.1005
R15661 a_21692_n6694.n7 a_21692_n6694.t9 16.3282
R15662 a_21692_n6694.n22 a_21692_n6694.t24 16.3282
R15663 a_21692_n6694.n4 a_21692_n6694.n2 15.8405
R15664 a_21692_n6694.n6 a_21692_n6694.t19 15.3305
R15665 a_21692_n6694.n6 a_21692_n6694.t15 15.148
R15666 a_21692_n6694.n13 a_21692_n6694.t35 14.7465
R15667 a_21692_n6694.n7 a_21692_n6694.t14 14.7465
R15668 a_21692_n6694.n22 a_21692_n6694.t33 14.7465
R15669 a_21692_n6694.n0 a_21692_n6694.n18 14.3221
R15670 a_21692_n6694.n15 a_21692_n6694.n11 12.7805
R15671 a_21692_n6694.n1 a_21692_n6694.n25 12.7371
R15672 a_21692_n6694.n28 a_21692_n6694.n27 12.6805
R15673 a_21692_n6694.n18 a_21692_n6694.t3 12.6782
R15674 a_21692_n6694.n23 a_21692_n6694.n22 12.5041
R15675 a_21692_n6694.n3 a_21692_n6694.t20 11.8873
R15676 a_21692_n6694.n25 a_21692_n6694.t2 11.8752
R15677 a_21692_n6694.n11 a_21692_n6694.n9 10.4405
R15678 a_21692_n6694.n0 a_21692_n6694.n17 10.0805
R15679 a_21692_n6694.n26 a_21692_n6694.n16 9.9005
R15680 a_21692_n6694.n0 a_21692_n6694.n19 9.9005
R15681 a_21692_n6694.n14 a_21692_n6694.n12 9.8129
R15682 a_21692_n6694.n9 a_21692_n6694.n8 9.4955
R15683 a_21692_n6694.n29 a_21692_n6694.n28 9.4055
R15684 a_21692_n6694.n4 a_21692_n6694.n3 8.58607
R15685 a_21692_n6694.n26 a_21692_n6694.n1 8.2805
R15686 a_21692_n6694.n14 a_21692_n6694.n13 8.0005
R15687 a_21692_n6694.n31 a_21692_n6694.t0 7.02633
R15688 a_21692_n6694.n16 a_21692_n6694.t10 6.71423
R15689 a_21692_n6694.n20 a_21692_n6694.t26 6.71423
R15690 a_21692_n6694.n17 a_21692_n6694.t32 6.71423
R15691 a_21692_n6694.n19 a_21692_n6694.t18 6.71423
R15692 a_21692_n6694.n2 a_21692_n6694.t12 6.71423
R15693 a_21692_n6694.n10 a_21692_n6694.t17 6.3005
R15694 a_21692_n6694.n5 a_21692_n6694.t8 6.3005
R15695 a_21692_n6694.n24 a_21692_n6694.t28 6.3005
R15696 a_21692_n6694.n30 a_21692_n6694.n29 6.3005
R15697 a_21692_n6694.n21 a_21692_n6694.n0 6.3005
R15698 a_21692_n6694.n29 a_21692_n6694.n15 5.9405
R15699 a_21692_n6694.n10 a_21692_n6694.t13 5.6196
R15700 a_21692_n6694.n5 a_21692_n6694.t6 5.6196
R15701 a_21692_n6694.n24 a_21692_n6694.t29 5.6196
R15702 a_21692_n6694.n28 a_21692_n6694.n26 5.5355
R15703 a_21692_n6694.n16 a_21692_n6694.t11 5.20587
R15704 a_21692_n6694.n20 a_21692_n6694.t23 5.20587
R15705 a_21692_n6694.n17 a_21692_n6694.t25 5.20587
R15706 a_21692_n6694.n19 a_21692_n6694.t21 5.20587
R15707 a_21692_n6694.n2 a_21692_n6694.t16 5.20587
R15708 a_21692_n6694.n15 a_21692_n6694.n14 4.58256
R15709 a_21692_n6694.n11 a_21692_n6694.n10 4.53811
R15710 a_21692_n6694.n9 a_21692_n6694.n5 4.53811
R15711 a_21692_n6694.n21 a_21692_n6694.n20 4.5005
R15712 a_21692_n6694.n31 a_21692_n6694.n30 4.5005
R15713 a_21692_n6694.n23 a_21692_n6694.n21 3.6455
R15714 a_21692_n6694.n1 a_21692_n6694.n23 2.8355
R15715 a_21692_n6694.t1 a_21692_n6694.n31 2.74964
R15716 a_24815_n3588.n11 a_24815_n3588.n10 26.1817
R15717 a_24815_n3588.n6 a_24815_n3588.t18 22.2655
R15718 a_24815_n3588.n9 a_24815_n3588.t5 18.6885
R15719 a_24815_n3588.n10 a_24815_n3588.t12 18.6155
R15720 a_24815_n3588.n15 a_24815_n3588.n12 17.9437
R15721 a_24815_n3588.n11 a_24815_n3588.n9 17.7217
R15722 a_24815_n3588.n12 a_24815_n3588.n8 17.5193
R15723 a_24815_n3588.n14 a_24815_n3588.t8 17.2772
R15724 a_24815_n3588.n7 a_24815_n3588.t13 16.5715
R15725 a_24815_n3588.n2 a_24815_n3588.n1 4.61819
R15726 a_24815_n3588.n14 a_24815_n3588.t9 16.4985
R15727 a_24815_n3588.n1 a_24815_n3588.t20 16.4985
R15728 a_24815_n3588.n3 a_24815_n3588.t15 16.4985
R15729 a_24815_n3588.n13 a_24815_n3588.t7 16.4985
R15730 a_24815_n3588.n13 a_24815_n3588.t14 15.6468
R15731 a_24815_n3588.n7 a_24815_n3588.t4 15.4643
R15732 a_24815_n3588.n8 a_24815_n3588.t17 15.3305
R15733 a_24815_n3588.n8 a_24815_n3588.t10 15.0872
R15734 a_24815_n3588.n0 a_24815_n3588.n5 14.9336
R15735 a_24815_n3588.n1 a_24815_n3588.t16 14.7952
R15736 a_24815_n3588.n3 a_24815_n3588.t19 14.7952
R15737 a_24815_n3588.n5 a_24815_n3588.t11 13.5573
R15738 a_24815_n3588.n9 a_24815_n3588.t6 11.8752
R15739 a_24815_n3588.n10 a_24815_n3588.t21 11.8752
R15740 a_24815_n3588.n16 a_24815_n3588.n0 11.6555
R15741 a_24815_n3588.n5 a_24815_n3588.t22 11.0235
R15742 a_24815_n3588.n2 a_24815_n3588.n3 4.61819
R15743 a_24815_n3588.n2 a_24815_n3588.n4 2.9334
R15744 a_24815_n3588.t3 a_24815_n3588.n16 9.9005
R15745 a_24815_n3588.t3 a_24815_n3588.t1 9.83456
R15746 a_24815_n3588.n6 a_24815_n3588.t23 9.77033
R15747 a_24815_n3588.n4 a_24815_n3588.n13 9.2005
R15748 a_24815_n3588.n16 a_24815_n3588.n15 9.1805
R15749 a_24815_n3588.n0 a_24815_n3588.n7 9.01391
R15750 a_24815_n3588.n12 a_24815_n3588.n11 8.6405
R15751 a_24815_n3588.n0 a_24815_n3588.n6 8.01708
R15752 a_24815_n3588.n4 a_24815_n3588.n14 8.0005
R15753 a_24815_n3588.t3 a_24815_n3588.t0 7.21149
R15754 a_24815_n3588.n15 a_24815_n3588.n4 6.25864
R15755 a_24815_n3588.t2 a_24815_n3588.t3 5.53329
R15756 a_45648_1564.n10 a_45648_1564.t10 15.8415
R15757 a_45648_1564.n4 a_45648_1564.t17 15.8415
R15758 a_45648_1564.n5 a_45648_1564.t9 15.8415
R15759 a_45648_1564.n6 a_45648_1564.t15 15.8415
R15760 a_45648_1564.n7 a_45648_1564.t16 15.8415
R15761 a_45648_1564.n8 a_45648_1564.t12 15.8415
R15762 a_45648_1564.n9 a_45648_1564.t13 15.8415
R15763 a_45648_1564.n11 a_45648_1564.t22 15.8415
R15764 a_45648_1564.n10 a_45648_1564.t20 13.4447
R15765 a_45648_1564.n4 a_45648_1564.t14 13.4447
R15766 a_45648_1564.n5 a_45648_1564.t19 13.4447
R15767 a_45648_1564.n6 a_45648_1564.t8 13.4447
R15768 a_45648_1564.n7 a_45648_1564.t11 13.4447
R15769 a_45648_1564.n8 a_45648_1564.t21 13.4447
R15770 a_45648_1564.n9 a_45648_1564.t23 13.4447
R15771 a_45648_1564.n11 a_45648_1564.t18 13.4447
R15772 a_45648_1564.n5 a_45648_1564.n4 10.5449
R15773 a_45648_1564.n6 a_45648_1564.n5 10.5449
R15774 a_45648_1564.n7 a_45648_1564.n6 10.5449
R15775 a_45648_1564.n8 a_45648_1564.n7 10.5449
R15776 a_45648_1564.n9 a_45648_1564.n8 10.5449
R15777 a_45648_1564.n11 a_45648_1564.n9 10.5449
R15778 a_45648_1564.n11 a_45648_1564.n10 10.5449
R15779 a_45648_1564.n0 a_45648_1564.n3 7.22489
R15780 a_45648_1564.n0 a_45648_1564.n2 6.36702
R15781 a_45648_1564.n12 a_45648_1564.n0 3.56115
R15782 a_45648_1564.n0 a_45648_1564.n1 2.68463
R15783 a_45648_1564.n0 a_45648_1564.n11 2.37315
R15784 a_45648_1564.n1 a_45648_1564.t6 2.06607
R15785 a_45648_1564.t7 a_45648_1564.n12 2.06607
R15786 a_45648_1564.n3 a_45648_1564.t0 1.99806
R15787 a_45648_1564.n3 a_45648_1564.t2 1.99806
R15788 a_45648_1564.n2 a_45648_1564.t3 1.99806
R15789 a_45648_1564.n2 a_45648_1564.t1 1.99806
R15790 a_45648_1564.n1 a_45648_1564.t4 1.4923
R15791 a_45648_1564.n12 a_45648_1564.t5 1.4923
R15792 EOC EOC.n14 9.97121
R15793 EOC.n11 EOC.n10 6.90733
R15794 EOC.n8 EOC.n7 6.89497
R15795 EOC.n11 EOC.n9 6.3768
R15796 EOC.n8 EOC.n6 6.3768
R15797 EOC.n2 EOC.n1 3.23472
R15798 EOC.n5 EOC.n4 3.21104
R15799 EOC.n5 EOC.n3 2.7042
R15800 EOC.n2 EOC.n0 2.7042
R15801 EOC.n3 EOC.t13 2.06607
R15802 EOC.n4 EOC.t14 2.06607
R15803 EOC.n1 EOC.t9 2.06607
R15804 EOC.n0 EOC.t11 2.06607
R15805 EOC.n9 EOC.t7 1.99806
R15806 EOC.n9 EOC.t6 1.99806
R15807 EOC.n10 EOC.t5 1.99806
R15808 EOC.n10 EOC.t3 1.99806
R15809 EOC.n7 EOC.t4 1.99806
R15810 EOC.n7 EOC.t2 1.99806
R15811 EOC.n6 EOC.t1 1.99806
R15812 EOC.n6 EOC.t0 1.99806
R15813 EOC.n3 EOC.t12 1.4923
R15814 EOC.n4 EOC.t8 1.4923
R15815 EOC.n1 EOC.t15 1.4923
R15816 EOC.n0 EOC.t10 1.4923
R15817 EOC.n12 EOC.n11 0.189974
R15818 EOC.n13 EOC.n5 0.175763
R15819 EOC.n12 EOC.n8 0.152079
R15820 EOC.n13 EOC.n12 0.145625
R15821 EOC.n14 EOC.n2 0.128395
R15822 EOC.n14 EOC.n13 0.0383947
R15823 a_22444_332.n0 a_22444_332.n4 30.9322
R15824 a_22444_332.t1 a_22444_332.n1 25.4705
R15825 a_22444_332.n14 a_22444_332.n13 22.9055
R15826 a_22444_332.t1 a_22444_332.n14 22.4105
R15827 a_22444_332.n0 a_22444_332.t11 20.9945
R15828 a_22444_332.n13 a_22444_332.n12 18.2821
R15829 a_22444_332.n6 a_22444_332.t29 17.7395
R15830 a_22444_332.n12 a_22444_332.t30 17.7395
R15831 a_22444_332.n9 a_22444_332.t23 17.7395
R15832 a_22444_332.n4 a_22444_332.t20 17.484
R15833 a_22444_332.n2 a_22444_332.t21 17.119
R15834 a_22444_332.n5 a_22444_332.t36 17.119
R15835 a_22444_332.n0 a_22444_332.t22 16.9182
R15836 a_22444_332.n7 a_22444_332.n6 16.6171
R15837 a_22444_332.n3 a_22444_332.t12 16.1822
R15838 a_22444_332.n3 a_22444_332.t32 14.0165
R15839 a_22444_332.n0 a_22444_332.n3 13.4207
R15840 a_22444_332.n10 a_22444_332.n9 13.0769
R15841 a_22444_332.n1 a_22444_332.n5 12.7446
R15842 a_22444_332.n2 a_22444_332.t8 12.7147
R15843 a_22444_332.n5 a_22444_332.t7 12.7147
R15844 a_22444_332.n6 a_22444_332.t13 12.6782
R15845 a_22444_332.n12 a_22444_332.t28 12.6782
R15846 a_22444_332.n9 a_22444_332.t17 12.6782
R15847 a_22444_332.n1 a_22444_332.n2 12.5914
R15848 a_22444_332.n4 a_22444_332.t14 11.863
R15849 a_22444_332.n7 a_22444_332.t27 11.6555
R15850 a_22444_332.t19 a_22444_332.t33 11.6038
R15851 a_22444_332.n1 a_22444_332.t19 11.2055
R15852 a_22444_332.t26 a_22444_332.t25 11.0638
R15853 a_22444_332.n1 a_22444_332.n8 10.9805
R15854 a_22444_332.n14 a_22444_332.n10 10.6537
R15855 a_22444_332.n8 a_22444_332.t26 9.7205
R15856 a_22444_332.n10 a_22444_332.t16 9.7205
R15857 a_22444_332.t19 a_22444_332.t15 9.3155
R15858 a_22444_332.t0 a_22444_332.t1 9.01572
R15859 a_22444_332.n8 a_22444_332.t10 9.0005
R15860 a_22444_332.t1 a_22444_332.t3 8.51574
R15861 a_22444_332.t19 a_22444_332.n0 8.4605
R15862 a_22444_332.t1 a_22444_332.t4 7.3492
R15863 a_22444_332.t27 a_22444_332.t31 6.71423
R15864 a_22444_332.t26 a_22444_332.n7 6.6605
R15865 a_22444_332.n13 a_22444_332.n11 6.65311
R15866 a_22444_332.t10 a_22444_332.t18 6.56378
R15867 a_22444_332.t15 a_22444_332.t34 6.41334
R15868 a_22444_332.t16 a_22444_332.t24 6.41334
R15869 a_22444_332.n11 a_22444_332.t9 6.3005
R15870 a_22444_332.t1 a_22444_332.t5 6.3005
R15871 a_22444_332.t1 a_22444_332.t6 6.07917
R15872 a_22444_332.t1 a_22444_332.t2 5.86452
R15873 a_22444_332.n11 a_22444_332.t35 5.6196
R15874 a_11087_n23528.n137 a_11087_n23528.n136 39.8544
R15875 a_11087_n23528.n1 a_11087_n23528.n2 0.47779
R15876 a_11087_n23528.n32 a_11087_n23528.n30 10.553
R15877 a_11087_n23528.n139 a_11087_n23528.n138 10.4369
R15878 a_11087_n23528.n141 a_11087_n23528.n140 10.4369
R15879 a_11087_n23528.n143 a_11087_n23528.n142 10.4308
R15880 a_11087_n23528.n145 a_11087_n23528.n144 10.4308
R15881 a_11087_n23528.n147 a_11087_n23528.n146 10.4308
R15882 a_11087_n23528.n32 a_11087_n23528.n31 10.4156
R15883 a_11087_n23528.n36 a_11087_n23528.n35 10.4129
R15884 a_11087_n23528.n38 a_11087_n23528.n37 10.4121
R15885 a_11087_n23528.n34 a_11087_n23528.n33 10.4121
R15886 a_11087_n23528.n23 a_11087_n23528.n21 10.357
R15887 a_11087_n23528.n29 a_11087_n23528.n28 10.2004
R15888 a_11087_n23528.n25 a_11087_n23528.n24 10.2004
R15889 a_11087_n23528.n27 a_11087_n23528.n26 10.198
R15890 a_11087_n23528.n23 a_11087_n23528.n22 10.1921
R15891 a_11087_n23528.n125 a_11087_n23528.n124 5.2655
R15892 a_11087_n23528.n131 a_11087_n23528.n90 4.5675
R15893 a_11087_n23528.n136 a_11087_n23528.n135 4.5675
R15894 a_11087_n23528.n130 a_11087_n23528.n129 4.5675
R15895 a_11087_n23528.n128 a_11087_n23528.n125 4.5675
R15896 a_11087_n23528.n101 a_11087_n23528.n2 3.39337
R15897 a_11087_n23528.n107 a_11087_n23528.n98 4.5675
R15898 a_11087_n23528.n112 a_11087_n23528.n111 4.5675
R15899 a_11087_n23528.n101 a_11087_n23528.n100 4.5675
R15900 a_11087_n23528.n106 a_11087_n23528.n105 4.5675
R15901 a_11087_n23528.n119 a_11087_n23528.n94 4.5675
R15902 a_11087_n23528.n124 a_11087_n23528.n123 4.5675
R15903 a_11087_n23528.n113 a_11087_n23528.n96 4.5675
R15904 a_11087_n23528.n118 a_11087_n23528.n117 4.5675
R15905 a_11087_n23528.n83 a_11087_n23528.n41 4.5675
R15906 a_11087_n23528.n77 a_11087_n23528.n43 4.5675
R15907 a_11087_n23528.n82 a_11087_n23528.n81 4.5675
R15908 a_11087_n23528.n88 a_11087_n23528.n87 4.5675
R15909 a_11087_n23528.n65 a_11087_n23528.n47 4.5675
R15910 a_11087_n23528.n70 a_11087_n23528.n69 4.5675
R15911 a_11087_n23528.n71 a_11087_n23528.n45 4.5675
R15912 a_11087_n23528.n76 a_11087_n23528.n75 4.5675
R15913 a_11087_n23528.n59 a_11087_n23528.n49 4.5675
R15914 a_11087_n23528.n64 a_11087_n23528.n63 4.5675
R15915 a_11087_n23528.n58 a_11087_n23528.n57 4.5675
R15916 a_11087_n23528.n55 a_11087_n23528.n52 4.5675
R15917 a_11087_n23528.n52 a_11087_n23528.t44 6.7695
R15918 a_11087_n23528.n103 a_11087_n23528.n102 4.5005
R15919 a_11087_n23528.n104 a_11087_n23528.n99 4.5005
R15920 a_11087_n23528.n109 a_11087_n23528.n108 4.5005
R15921 a_11087_n23528.n110 a_11087_n23528.n97 4.5005
R15922 a_11087_n23528.n115 a_11087_n23528.n114 4.5005
R15923 a_11087_n23528.n116 a_11087_n23528.n95 4.5005
R15924 a_11087_n23528.n121 a_11087_n23528.n120 4.5005
R15925 a_11087_n23528.n122 a_11087_n23528.n93 4.5005
R15926 a_11087_n23528.n127 a_11087_n23528.n126 4.5005
R15927 a_11087_n23528.n92 a_11087_n23528.n91 4.5005
R15928 a_11087_n23528.n133 a_11087_n23528.n132 4.5005
R15929 a_11087_n23528.n134 a_11087_n23528.n89 4.5005
R15930 a_11087_n23528.n54 a_11087_n23528.n53 4.5005
R15931 a_11087_n23528.n51 a_11087_n23528.n50 4.5005
R15932 a_11087_n23528.n61 a_11087_n23528.n60 4.5005
R15933 a_11087_n23528.n62 a_11087_n23528.n48 4.5005
R15934 a_11087_n23528.n67 a_11087_n23528.n66 4.5005
R15935 a_11087_n23528.n68 a_11087_n23528.n46 4.5005
R15936 a_11087_n23528.n73 a_11087_n23528.n72 4.5005
R15937 a_11087_n23528.n74 a_11087_n23528.n44 4.5005
R15938 a_11087_n23528.n79 a_11087_n23528.n78 4.5005
R15939 a_11087_n23528.n80 a_11087_n23528.n42 4.5005
R15940 a_11087_n23528.n85 a_11087_n23528.n84 4.5005
R15941 a_11087_n23528.n86 a_11087_n23528.n40 4.5005
R15942 a_11087_n23528.n135 a_11087_n23528.n5 2.21775
R15943 a_11087_n23528.n90 a_11087_n23528.n5 2.21775
R15944 a_11087_n23528.t50 a_11087_n23528.n128 2.21775
R15945 a_11087_n23528.n129 a_11087_n23528.t50 2.21775
R15946 a_11087_n23528.n111 a_11087_n23528.n1 2.21775
R15947 a_11087_n23528.n98 a_11087_n23528.n1 2.21775
R15948 a_11087_n23528.n105 a_11087_n23528.n1 2.21775
R15949 a_11087_n23528.n100 a_11087_n23528.n1 2.21775
R15950 a_11087_n23528.n123 a_11087_n23528.n18 2.21775
R15951 a_11087_n23528.n94 a_11087_n23528.n18 2.21775
R15952 a_11087_n23528.n117 a_11087_n23528.n19 2.21775
R15953 a_11087_n23528.n96 a_11087_n23528.n19 2.21775
R15954 a_11087_n23528.n81 a_11087_n23528.t35 2.21775
R15955 a_11087_n23528.n43 a_11087_n23528.t35 2.21775
R15956 a_11087_n23528.n87 a_11087_n23528.t35 2.21775
R15957 a_11087_n23528.n41 a_11087_n23528.t35 2.21775
R15958 a_11087_n23528.n69 a_11087_n23528.n0 2.21775
R15959 a_11087_n23528.n47 a_11087_n23528.n0 2.21775
R15960 a_11087_n23528.n75 a_11087_n23528.n0 2.21775
R15961 a_11087_n23528.n45 a_11087_n23528.n0 2.21775
R15962 a_11087_n23528.n63 a_11087_n23528.n16 2.21775
R15963 a_11087_n23528.n49 a_11087_n23528.n16 2.21775
R15964 a_11087_n23528.n56 a_11087_n23528.n55 2.21775
R15965 a_11087_n23528.n57 a_11087_n23528.n56 2.21775
R15966 a_11087_n23528.n113 a_11087_n23528.n112 1.8905
R15967 a_11087_n23528.n77 a_11087_n23528.n76 1.8905
R15968 a_11087_n23528.n65 a_11087_n23528.n64 1.88938
R15969 a_11087_n23528.n137 a_11087_n23528.n88 1.68967
R15970 a_11087_n23528.n139 a_11087_n23528.n137 1.51044
R15971 a_11087_n23528.n15 a_11087_n23528.n6 0.0144139
R15972 a_11087_n23528.n6 a_11087_n23528.t43 0.495679
R15973 a_11087_n23528.t50 a_11087_n23528.n3 0.471104
R15974 a_11087_n23528.n10 a_11087_n23528.n9 0.0280721
R15975 a_11087_n23528.n9 a_11087_n23528.t31 0.467713
R15976 a_11087_n23528.n4 a_11087_n23528.t38 0.474486
R15977 a_11087_n23528.n3 a_11087_n23528.n4 0.0274329
R15978 a_11087_n23528.n7 a_11087_n23528.t59 0.467464
R15979 a_11087_n23528.n8 a_11087_n23528.n7 0.0280716
R15980 a_11087_n23528.n13 a_11087_n23528.n14 0.0280716
R15981 a_11087_n23528.n14 a_11087_n23528.t55 0.467464
R15982 a_11087_n23528.n11 a_11087_n23528.n12 0.0280716
R15983 a_11087_n23528.n12 a_11087_n23528.t37 0.467464
R15984 a_11087_n23528.n39 a_11087_n23528.n29 0.773592
R15985 a_11087_n23528.n107 a_11087_n23528.n106 0.676625
R15986 a_11087_n23528.n59 a_11087_n23528.n58 0.676625
R15987 a_11087_n23528.n131 a_11087_n23528.n130 0.6755
R15988 a_11087_n23528.n119 a_11087_n23528.n118 0.6755
R15989 a_11087_n23528.n83 a_11087_n23528.n82 0.6755
R15990 a_11087_n23528.n71 a_11087_n23528.n70 0.6755
R15991 a_11087_n23528.n28 a_11087_n23528.t12 0.6505
R15992 a_11087_n23528.n28 a_11087_n23528.t16 0.6505
R15993 a_11087_n23528.n26 a_11087_n23528.t11 0.6505
R15994 a_11087_n23528.n26 a_11087_n23528.t19 0.6505
R15995 a_11087_n23528.n24 a_11087_n23528.t14 0.6505
R15996 a_11087_n23528.n24 a_11087_n23528.t18 0.6505
R15997 a_11087_n23528.n22 a_11087_n23528.t17 0.6505
R15998 a_11087_n23528.n22 a_11087_n23528.t10 0.6505
R15999 a_11087_n23528.n21 a_11087_n23528.t15 0.6505
R16000 a_11087_n23528.n21 a_11087_n23528.t13 0.6505
R16001 a_11087_n23528.t54 a_11087_n23528.t34 0.610813
R16002 a_11087_n23528.t58 a_11087_n23528.t61 0.610813
R16003 a_11087_n23528.n138 a_11087_n23528.t21 0.5855
R16004 a_11087_n23528.n138 a_11087_n23528.t25 0.5855
R16005 a_11087_n23528.n140 a_11087_n23528.t24 0.5855
R16006 a_11087_n23528.n140 a_11087_n23528.t28 0.5855
R16007 a_11087_n23528.n142 a_11087_n23528.t27 0.5855
R16008 a_11087_n23528.n142 a_11087_n23528.t20 0.5855
R16009 a_11087_n23528.n144 a_11087_n23528.t26 0.5855
R16010 a_11087_n23528.n144 a_11087_n23528.t23 0.5855
R16011 a_11087_n23528.n37 a_11087_n23528.t9 0.5855
R16012 a_11087_n23528.n37 a_11087_n23528.t3 0.5855
R16013 a_11087_n23528.n35 a_11087_n23528.t8 0.5855
R16014 a_11087_n23528.n35 a_11087_n23528.t6 0.5855
R16015 a_11087_n23528.n33 a_11087_n23528.t1 0.5855
R16016 a_11087_n23528.n33 a_11087_n23528.t5 0.5855
R16017 a_11087_n23528.n31 a_11087_n23528.t4 0.5855
R16018 a_11087_n23528.n31 a_11087_n23528.t7 0.5855
R16019 a_11087_n23528.n30 a_11087_n23528.t2 0.5855
R16020 a_11087_n23528.n30 a_11087_n23528.t0 0.5855
R16021 a_11087_n23528.t29 a_11087_n23528.n147 0.5855
R16022 a_11087_n23528.n147 a_11087_n23528.t22 0.5855
R16023 a_11087_n23528.t53 a_11087_n23528.t42 0.582955
R16024 a_11087_n23528.n8 a_11087_n23528.t40 0.582955
R16025 a_11087_n23528.n12 a_11087_n23528.t41 0.610527
R16026 a_11087_n23528.t44 a_11087_n23528.n6 0.581013
R16027 a_11087_n23528.n0 a_11087_n23528.t35 0.550768
R16028 a_11087_n23528.t36 a_11087_n23528.t51 0.5405
R16029 a_11087_n23528.t33 a_11087_n23528.t46 0.5405
R16030 a_11087_n23528.n4 a_11087_n23528.t54 0.540346
R16031 a_11087_n23528.n10 a_11087_n23528.t36 0.512643
R16032 a_11087_n23528.n14 a_11087_n23528.t33 0.540214
R16033 a_11087_n23528.n15 a_11087_n23528.t58 0.512643
R16034 a_11087_n23528.t51 a_11087_n23528.n7 0.540214
R16035 a_11087_n23528.t46 a_11087_n23528.n11 0.512643
R16036 a_11087_n23528.n1 a_11087_n23528.n20 0.501102
R16037 a_11087_n23528.n17 a_11087_n23528.n0 0.499684
R16038 a_11087_n23528.t35 a_11087_n23528.n13 0.513368
R16039 a_11087_n23528.n39 a_11087_n23528.n38 0.366893
R16040 a_11087_n23528.n146 a_11087_n23528.n39 0.297718
R16041 a_11087_n23528.n141 a_11087_n23528.n139 0.1615
R16042 a_11087_n23528.n29 a_11087_n23528.n27 0.161
R16043 a_11087_n23528.n25 a_11087_n23528.n23 0.1605
R16044 a_11087_n23528.n27 a_11087_n23528.n25 0.1605
R16045 a_11087_n23528.n146 a_11087_n23528.n145 0.1605
R16046 a_11087_n23528.n145 a_11087_n23528.n143 0.1605
R16047 a_11087_n23528.n143 a_11087_n23528.n141 0.1585
R16048 a_11087_n23528.n38 a_11087_n23528.n36 0.139126
R16049 a_11087_n23528.n34 a_11087_n23528.n32 0.136566
R16050 a_11087_n23528.n134 a_11087_n23528.n133 0.1355
R16051 a_11087_n23528.n127 a_11087_n23528.n92 0.1355
R16052 a_11087_n23528.n110 a_11087_n23528.n109 0.1355
R16053 a_11087_n23528.n104 a_11087_n23528.n103 0.1355
R16054 a_11087_n23528.n122 a_11087_n23528.n121 0.1355
R16055 a_11087_n23528.n116 a_11087_n23528.n115 0.1355
R16056 a_11087_n23528.n136 a_11087_n23528.n89 0.1355
R16057 a_11087_n23528.n132 a_11087_n23528.n89 0.1355
R16058 a_11087_n23528.n132 a_11087_n23528.n131 0.1355
R16059 a_11087_n23528.n130 a_11087_n23528.n91 0.1355
R16060 a_11087_n23528.n126 a_11087_n23528.n91 0.1355
R16061 a_11087_n23528.n126 a_11087_n23528.n125 0.1355
R16062 a_11087_n23528.n124 a_11087_n23528.n93 0.1355
R16063 a_11087_n23528.n120 a_11087_n23528.n93 0.1355
R16064 a_11087_n23528.n120 a_11087_n23528.n119 0.1355
R16065 a_11087_n23528.n118 a_11087_n23528.n95 0.1355
R16066 a_11087_n23528.n114 a_11087_n23528.n95 0.1355
R16067 a_11087_n23528.n114 a_11087_n23528.n113 0.1355
R16068 a_11087_n23528.n112 a_11087_n23528.n97 0.1355
R16069 a_11087_n23528.n108 a_11087_n23528.n97 0.1355
R16070 a_11087_n23528.n108 a_11087_n23528.n107 0.1355
R16071 a_11087_n23528.n106 a_11087_n23528.n99 0.1355
R16072 a_11087_n23528.n102 a_11087_n23528.n99 0.1355
R16073 a_11087_n23528.n102 a_11087_n23528.n101 0.1355
R16074 a_11087_n23528.n86 a_11087_n23528.n85 0.1355
R16075 a_11087_n23528.n80 a_11087_n23528.n79 0.1355
R16076 a_11087_n23528.n68 a_11087_n23528.n67 0.1355
R16077 a_11087_n23528.n74 a_11087_n23528.n73 0.1355
R16078 a_11087_n23528.n62 a_11087_n23528.n61 0.1355
R16079 a_11087_n23528.n54 a_11087_n23528.n51 0.1355
R16080 a_11087_n23528.n88 a_11087_n23528.n40 0.1355
R16081 a_11087_n23528.n84 a_11087_n23528.n40 0.1355
R16082 a_11087_n23528.n84 a_11087_n23528.n83 0.1355
R16083 a_11087_n23528.n82 a_11087_n23528.n42 0.1355
R16084 a_11087_n23528.n78 a_11087_n23528.n42 0.1355
R16085 a_11087_n23528.n78 a_11087_n23528.n77 0.1355
R16086 a_11087_n23528.n76 a_11087_n23528.n44 0.1355
R16087 a_11087_n23528.n72 a_11087_n23528.n44 0.1355
R16088 a_11087_n23528.n72 a_11087_n23528.n71 0.1355
R16089 a_11087_n23528.n70 a_11087_n23528.n46 0.1355
R16090 a_11087_n23528.n66 a_11087_n23528.n46 0.1355
R16091 a_11087_n23528.n66 a_11087_n23528.n65 0.1355
R16092 a_11087_n23528.n64 a_11087_n23528.n48 0.1355
R16093 a_11087_n23528.n60 a_11087_n23528.n48 0.1355
R16094 a_11087_n23528.n60 a_11087_n23528.n59 0.1355
R16095 a_11087_n23528.n58 a_11087_n23528.n50 0.1355
R16096 a_11087_n23528.n53 a_11087_n23528.n50 0.1355
R16097 a_11087_n23528.n53 a_11087_n23528.n52 0.1355
R16098 a_11087_n23528.n36 a_11087_n23528.n34 0.13486
R16099 a_11087_n23528.n17 a_11087_n23528.n16 0.0773679
R16100 a_11087_n23528.n20 a_11087_n23528.n18 0.0762987
R16101 a_11087_n23528.n56 a_11087_n23528.n17 0.0762987
R16102 a_11087_n23528.n20 a_11087_n23528.n19 0.0762987
R16103 a_11087_n23528.n3 a_11087_n23528.t49 0.0708125
R16104 a_11087_n23528.n20 a_11087_n23528.t45 0.0708125
R16105 a_11087_n23528.n8 a_11087_n23528.t52 0.0708125
R16106 a_11087_n23528.n10 a_11087_n23528.t48 0.0708125
R16107 a_11087_n23528.n11 a_11087_n23528.t56 0.0708125
R16108 a_11087_n23528.n13 a_11087_n23528.t47 0.0708125
R16109 a_11087_n23528.n17 a_11087_n23528.t32 0.0708125
R16110 a_11087_n23528.n15 a_11087_n23528.t30 0.0708125
R16111 a_11087_n23528.n135 a_11087_n23528.n134 0.0675025
R16112 a_11087_n23528.n133 a_11087_n23528.n90 0.0675025
R16113 a_11087_n23528.n129 a_11087_n23528.n92 0.0675025
R16114 a_11087_n23528.n128 a_11087_n23528.n127 0.0675025
R16115 a_11087_n23528.n111 a_11087_n23528.n110 0.0675025
R16116 a_11087_n23528.n109 a_11087_n23528.n98 0.0675025
R16117 a_11087_n23528.n105 a_11087_n23528.n104 0.0675025
R16118 a_11087_n23528.n103 a_11087_n23528.n100 0.0675025
R16119 a_11087_n23528.n123 a_11087_n23528.n122 0.0675025
R16120 a_11087_n23528.n121 a_11087_n23528.n94 0.0675025
R16121 a_11087_n23528.n117 a_11087_n23528.n116 0.0675025
R16122 a_11087_n23528.n115 a_11087_n23528.n96 0.0675025
R16123 a_11087_n23528.n87 a_11087_n23528.n86 0.0675025
R16124 a_11087_n23528.n81 a_11087_n23528.n80 0.0675025
R16125 a_11087_n23528.n79 a_11087_n23528.n43 0.0675025
R16126 a_11087_n23528.n85 a_11087_n23528.n41 0.0675025
R16127 a_11087_n23528.n69 a_11087_n23528.n68 0.0675025
R16128 a_11087_n23528.n67 a_11087_n23528.n47 0.0675025
R16129 a_11087_n23528.n75 a_11087_n23528.n74 0.0675025
R16130 a_11087_n23528.n73 a_11087_n23528.n45 0.0675025
R16131 a_11087_n23528.n63 a_11087_n23528.n62 0.0675025
R16132 a_11087_n23528.n61 a_11087_n23528.n49 0.0675025
R16133 a_11087_n23528.n57 a_11087_n23528.n51 0.0675025
R16134 a_11087_n23528.n55 a_11087_n23528.n54 0.0675025
R16135 a_11087_n23528.n2 a_11087_n23528.n9 0.540956
R16136 a_11087_n23528.t53 a_11087_n23528.t38 0.501521
R16137 a_11087_n23528.n0 a_11087_n23528.t39 0.231838
R16138 a_11087_n23528.n1 a_11087_n23528.t60 0.223522
R16139 a_11087_n23528.n2 a_11087_n23528.t57 0.154606
R16140 a_11087_n23528.t50 a_11087_n23528.n5 0.152097
R16141 a_2167_3472.n9 a_2167_3472.t84 61.5517
R16142 a_2167_3472.n0 a_2167_3472.t1 15.8618
R16143 a_2167_3472.n0 a_2167_3472.t8 15.8393
R16144 a_2167_3472.n0 a_2167_3472.t32 15.7535
R16145 a_2167_3472.n0 a_2167_3472.t39 15.7496
R16146 a_2167_3472.n0 a_2167_3472.n1 14.963
R16147 a_2167_3472.n0 a_2167_3472.n3 14.9583
R16148 a_2167_3472.n0 a_2167_3472.n7 14.9559
R16149 a_2167_3472.n0 a_2167_3472.n6 14.9547
R16150 a_2167_3472.n0 a_2167_3472.n2 14.7096
R16151 a_2167_3472.n0 a_2167_3472.n5 14.7035
R16152 a_2167_3472.n0 a_2167_3472.n4 14.7035
R16153 a_2167_3472.n0 a_2167_3472.n8 14.6941
R16154 a_2167_3472.n9 a_2167_3472.n0 3.73147
R16155 a_2167_3472.t19 a_2167_3472.n9 3.13216
R16156 a_2167_3472.t19 a_2167_3472.t18 1.23983
R16157 a_2167_3472.t18 a_2167_3472.t24 1.23983
R16158 a_2167_3472.t24 a_2167_3472.t52 1.23983
R16159 a_2167_3472.t45 a_2167_3472.t42 1.23983
R16160 a_2167_3472.t42 a_2167_3472.t57 1.23983
R16161 a_2167_3472.t46 a_2167_3472.t65 1.23216
R16162 a_2167_3472.t63 a_2167_3472.t70 1.23216
R16163 a_2167_3472.t70 a_2167_3472.t27 1.23216
R16164 a_2167_3472.t80 a_2167_3472.t16 1.23216
R16165 a_2167_3472.t17 a_2167_3472.t12 1.23216
R16166 a_2167_3472.t26 a_2167_3472.t30 1.23216
R16167 a_2167_3472.t81 a_2167_3472.t49 1.23216
R16168 a_2167_3472.t78 a_2167_3472.t64 1.23216
R16169 a_2167_3472.t48 a_2167_3472.t53 1.23216
R16170 a_2167_3472.t48 a_2167_3472.t68 1.23216
R16171 a_2167_3472.t68 a_2167_3472.t74 1.23216
R16172 a_2167_3472.t52 a_2167_3472.t28 1.23216
R16173 a_2167_3472.t71 a_2167_3472.t29 1.23216
R16174 a_2167_3472.t75 a_2167_3472.t23 1.23216
R16175 a_2167_3472.t14 a_2167_3472.t15 1.23216
R16176 a_2167_3472.t83 a_2167_3472.t43 1.23216
R16177 a_2167_3472.t21 a_2167_3472.t58 1.23216
R16178 a_2167_3472.t72 a_2167_3472.t44 1.23216
R16179 a_2167_3472.t22 a_2167_3472.t21 1.23216
R16180 a_2167_3472.t22 a_2167_3472.t20 1.23216
R16181 a_2167_3472.t73 a_2167_3472.t41 1.23216
R16182 a_2167_3472.t62 a_2167_3472.t13 1.23216
R16183 a_2167_3472.t43 a_2167_3472.t50 1.23216
R16184 a_2167_3472.t14 a_2167_3472.t51 1.23216
R16185 a_2167_3472.t75 a_2167_3472.t66 1.23216
R16186 a_2167_3472.t71 a_2167_3472.t54 1.23216
R16187 a_2167_3472.t28 a_2167_3472.t57 1.23216
R16188 a_2167_3472.t30 a_2167_3472.t12 1.2245
R16189 a_2167_3472.t83 a_2167_3472.t76 1.2245
R16190 a_2167_3472.t49 a_2167_3472.t30 1.2245
R16191 a_2167_3472.t83 a_2167_3472.t15 1.2245
R16192 a_2167_3472.t64 a_2167_3472.t49 1.2245
R16193 a_2167_3472.t15 a_2167_3472.t23 1.2245
R16194 a_2167_3472.t53 a_2167_3472.t64 1.2245
R16195 a_2167_3472.t23 a_2167_3472.t29 1.2245
R16196 a_2167_3472.t52 a_2167_3472.t53 1.2245
R16197 a_2167_3472.t61 a_2167_3472.t11 1.2245
R16198 a_2167_3472.t55 a_2167_3472.t67 1.2245
R16199 a_2167_3472.t69 a_2167_3472.t55 1.2245
R16200 a_2167_3472.t56 a_2167_3472.t69 1.2245
R16201 a_2167_3472.t61 a_2167_3472.t46 1.2245
R16202 a_2167_3472.t46 a_2167_3472.t56 1.2245
R16203 a_2167_3472.t11 a_2167_3472.t65 1.2245
R16204 a_2167_3472.t65 a_2167_3472.t25 1.2245
R16205 a_2167_3472.t56 a_2167_3472.t25 1.2245
R16206 a_2167_3472.t25 a_2167_3472.t79 1.2245
R16207 a_2167_3472.t69 a_2167_3472.t79 1.2245
R16208 a_2167_3472.t79 a_2167_3472.t47 1.2245
R16209 a_2167_3472.t55 a_2167_3472.t47 1.2245
R16210 a_2167_3472.t63 a_2167_3472.t47 1.2245
R16211 a_2167_3472.t67 a_2167_3472.t63 1.2245
R16212 a_2167_3472.t27 a_2167_3472.t58 1.2245
R16213 a_2167_3472.t72 a_2167_3472.t80 1.2245
R16214 a_2167_3472.t80 a_2167_3472.t27 1.2245
R16215 a_2167_3472.t80 a_2167_3472.t12 1.2245
R16216 a_2167_3472.t16 a_2167_3472.t70 1.2245
R16217 a_2167_3472.t16 a_2167_3472.t47 1.2245
R16218 a_2167_3472.t16 a_2167_3472.t17 1.2245
R16219 a_2167_3472.t17 a_2167_3472.t79 1.2245
R16220 a_2167_3472.t17 a_2167_3472.t26 1.2245
R16221 a_2167_3472.t26 a_2167_3472.t25 1.2245
R16222 a_2167_3472.t26 a_2167_3472.t81 1.2245
R16223 a_2167_3472.t81 a_2167_3472.t65 1.2245
R16224 a_2167_3472.t81 a_2167_3472.t78 1.2245
R16225 a_2167_3472.t78 a_2167_3472.t11 1.2245
R16226 a_2167_3472.t78 a_2167_3472.t48 1.2245
R16227 a_2167_3472.t48 a_2167_3472.t24 1.2245
R16228 a_2167_3472.t68 a_2167_3472.t11 1.2245
R16229 a_2167_3472.t68 a_2167_3472.t18 1.2245
R16230 a_2167_3472.t74 a_2167_3472.t61 1.2245
R16231 a_2167_3472.t74 a_2167_3472.t19 1.2245
R16232 a_2167_3472.t29 a_2167_3472.t57 1.2245
R16233 a_2167_3472.t76 a_2167_3472.t44 1.2245
R16234 a_2167_3472.t21 a_2167_3472.t44 1.2245
R16235 a_2167_3472.t73 a_2167_3472.t20 1.2245
R16236 a_2167_3472.t41 a_2167_3472.t22 1.2245
R16237 a_2167_3472.t41 a_2167_3472.t44 1.2245
R16238 a_2167_3472.t43 a_2167_3472.t13 1.2245
R16239 a_2167_3472.t41 a_2167_3472.t13 1.2245
R16240 a_2167_3472.t13 a_2167_3472.t76 1.2245
R16241 a_2167_3472.t62 a_2167_3472.t73 1.2245
R16242 a_2167_3472.t50 a_2167_3472.t62 1.2245
R16243 a_2167_3472.t66 a_2167_3472.t51 1.2245
R16244 a_2167_3472.t51 a_2167_3472.t50 1.2245
R16245 a_2167_3472.t43 a_2167_3472.t14 1.2245
R16246 a_2167_3472.t14 a_2167_3472.t75 1.2245
R16247 a_2167_3472.t71 a_2167_3472.t42 1.2245
R16248 a_2167_3472.t75 a_2167_3472.t71 1.2245
R16249 a_2167_3472.t54 a_2167_3472.t66 1.2245
R16250 a_2167_3472.t54 a_2167_3472.t45 1.2245
R16251 a_2167_3472.t28 a_2167_3472.t77 1.2245
R16252 a_2167_3472.t77 a_2167_3472.t29 1.2245
R16253 a_2167_3472.t77 a_2167_3472.t53 1.2245
R16254 a_2167_3472.t77 a_2167_3472.t10 1.2245
R16255 a_2167_3472.t10 a_2167_3472.t23 1.2245
R16256 a_2167_3472.t10 a_2167_3472.t64 1.2245
R16257 a_2167_3472.t10 a_2167_3472.t60 1.2245
R16258 a_2167_3472.t60 a_2167_3472.t15 1.2245
R16259 a_2167_3472.t60 a_2167_3472.t49 1.2245
R16260 a_2167_3472.t60 a_2167_3472.t82 1.2245
R16261 a_2167_3472.t82 a_2167_3472.t83 1.2245
R16262 a_2167_3472.t82 a_2167_3472.t30 1.2245
R16263 a_2167_3472.t82 a_2167_3472.t59 1.2245
R16264 a_2167_3472.t76 a_2167_3472.t59 1.2245
R16265 a_2167_3472.t12 a_2167_3472.t59 1.2245
R16266 a_2167_3472.t72 a_2167_3472.t59 1.2245
R16267 a_2167_3472.t72 a_2167_3472.t58 1.2245
R16268 a_2167_3472.n8 a_2167_3472.t35 0.6505
R16269 a_2167_3472.n8 a_2167_3472.t38 0.6505
R16270 a_2167_3472.n5 a_2167_3472.t36 0.6505
R16271 a_2167_3472.n5 a_2167_3472.t31 0.6505
R16272 a_2167_3472.n4 a_2167_3472.t40 0.6505
R16273 a_2167_3472.n4 a_2167_3472.t33 0.6505
R16274 a_2167_3472.n2 a_2167_3472.t34 0.6505
R16275 a_2167_3472.n2 a_2167_3472.t37 0.6505
R16276 a_2167_3472.n7 a_2167_3472.t4 0.5855
R16277 a_2167_3472.n7 a_2167_3472.t7 0.5855
R16278 a_2167_3472.n6 a_2167_3472.t5 0.5855
R16279 a_2167_3472.n6 a_2167_3472.t0 0.5855
R16280 a_2167_3472.n3 a_2167_3472.t9 0.5855
R16281 a_2167_3472.n3 a_2167_3472.t2 0.5855
R16282 a_2167_3472.n1 a_2167_3472.t3 0.5855
R16283 a_2167_3472.n1 a_2167_3472.t6 0.5855
R16284 a_21772_1116.n2 a_21772_1116.t17 15.8415
R16285 a_21772_1116.n3 a_21772_1116.t16 15.8415
R16286 a_21772_1116.n4 a_21772_1116.t4 15.8415
R16287 a_21772_1116.n5 a_21772_1116.t18 15.8415
R16288 a_21772_1116.n6 a_21772_1116.t15 15.8415
R16289 a_21772_1116.n7 a_21772_1116.t14 15.8415
R16290 a_21772_1116.n1 a_21772_1116.t5 15.8415
R16291 a_21772_1116.n0 a_21772_1116.t19 15.8415
R16292 a_21772_1116.n2 a_21772_1116.t8 13.4447
R16293 a_21772_1116.n3 a_21772_1116.t6 13.4447
R16294 a_21772_1116.n4 a_21772_1116.t12 13.4447
R16295 a_21772_1116.n5 a_21772_1116.t9 13.4447
R16296 a_21772_1116.n6 a_21772_1116.t7 13.4447
R16297 a_21772_1116.n7 a_21772_1116.t11 13.4447
R16298 a_21772_1116.n1 a_21772_1116.t13 13.4447
R16299 a_21772_1116.n0 a_21772_1116.t10 13.4447
R16300 a_21772_1116.n3 a_21772_1116.n2 10.5449
R16301 a_21772_1116.n4 a_21772_1116.n3 10.5449
R16302 a_21772_1116.n5 a_21772_1116.n4 10.5449
R16303 a_21772_1116.n6 a_21772_1116.n5 10.5449
R16304 a_21772_1116.n7 a_21772_1116.n6 10.5449
R16305 a_21772_1116.n0 a_21772_1116.n1 10.5449
R16306 a_21772_1116.n0 a_21772_1116.n7 10.5449
R16307 a_21772_1116.n0 a_21772_1116.t2 7.22489
R16308 a_21772_1116.n0 a_21772_1116.t3 7.12153
R16309 a_21772_1116.n0 a_21772_1116.t1 6.36702
R16310 a_21772_1116.t0 a_21772_1116.n0 5.62673
R16311 a_13623_n4162.n0 a_13623_n4162.t35 56.1018
R16312 a_13623_n4162.n1 a_13623_n4162.t22 56.0719
R16313 a_13623_n4162.n0 a_13623_n4162.t30 56.0141
R16314 a_13623_n4162.n0 a_13623_n4162.t27 55.9719
R16315 a_13623_n4162.n0 a_13623_n4162.t45 55.9719
R16316 a_13623_n4162.n0 a_13623_n4162.t37 55.9719
R16317 a_13623_n4162.n0 a_13623_n4162.t20 55.9719
R16318 a_13623_n4162.n0 a_13623_n4162.t42 55.9719
R16319 a_13623_n4162.n0 a_13623_n4162.t33 55.9719
R16320 a_13623_n4162.n0 a_13623_n4162.t18 55.9719
R16321 a_13623_n4162.n0 a_13623_n4162.t44 55.9719
R16322 a_13623_n4162.n0 a_13623_n4162.t23 55.9719
R16323 a_13623_n4162.n0 a_13623_n4162.t24 55.9719
R16324 a_13623_n4162.n0 a_13623_n4162.t41 55.9719
R16325 a_13623_n4162.n0 a_13623_n4162.t32 55.9719
R16326 a_13623_n4162.n0 a_13623_n4162.t17 55.9719
R16327 a_13623_n4162.n0 a_13623_n4162.t38 55.9719
R16328 a_13623_n4162.n0 a_13623_n4162.t29 55.9719
R16329 a_13623_n4162.n0 a_13623_n4162.t16 55.9719
R16330 a_13623_n4162.n0 a_13623_n4162.t40 55.9719
R16331 a_13623_n4162.n0 a_13623_n4162.t21 55.9719
R16332 a_13623_n4162.n1 a_13623_n4162.t36 55.9719
R16333 a_13623_n4162.n1 a_13623_n4162.t28 55.9719
R16334 a_13623_n4162.n1 a_13623_n4162.t19 55.9719
R16335 a_13623_n4162.n1 a_13623_n4162.t31 55.9719
R16336 a_13623_n4162.n1 a_13623_n4162.t25 55.9719
R16337 a_13623_n4162.n1 a_13623_n4162.t43 55.9719
R16338 a_13623_n4162.n4 a_13623_n4162.t34 55.9719
R16339 a_13623_n4162.n4 a_13623_n4162.t26 55.9719
R16340 a_13623_n4162.n4 a_13623_n4162.t39 55.9719
R16341 a_13623_n4162.n12 a_13623_n4162.n0 36.9047
R16342 a_13623_n4162.n3 a_13623_n4162.n8 6.90733
R16343 a_13623_n4162.n2 a_13623_n4162.n10 6.89497
R16344 a_13623_n4162.n2 a_13623_n4162.n9 6.3768
R16345 a_13623_n4162.n3 a_13623_n4162.n7 6.3768
R16346 a_13623_n4162.n3 a_13623_n4162.n6 3.21104
R16347 a_13623_n4162.n3 a_13623_n4162.n5 2.7042
R16348 a_13623_n4162.n13 a_13623_n4162.n3 2.7042
R16349 a_13623_n4162.n12 a_13623_n4162.n11 2.6005
R16350 a_13623_n4162.n6 a_13623_n4162.t14 2.06607
R16351 a_13623_n4162.n5 a_13623_n4162.t12 2.06607
R16352 a_13623_n4162.n11 a_13623_n4162.t10 2.06607
R16353 a_13623_n4162.t15 a_13623_n4162.n13 2.06607
R16354 a_13623_n4162.n9 a_13623_n4162.t2 1.99806
R16355 a_13623_n4162.n9 a_13623_n4162.t6 1.99806
R16356 a_13623_n4162.n10 a_13623_n4162.t0 1.99806
R16357 a_13623_n4162.n10 a_13623_n4162.t3 1.99806
R16358 a_13623_n4162.n8 a_13623_n4162.t7 1.99806
R16359 a_13623_n4162.n8 a_13623_n4162.t5 1.99806
R16360 a_13623_n4162.n7 a_13623_n4162.t4 1.99806
R16361 a_13623_n4162.n7 a_13623_n4162.t1 1.99806
R16362 a_13623_n4162.n6 a_13623_n4162.t8 1.4923
R16363 a_13623_n4162.n5 a_13623_n4162.t13 1.4923
R16364 a_13623_n4162.n11 a_13623_n4162.t11 1.4923
R16365 a_13623_n4162.n13 a_13623_n4162.t9 1.4923
R16366 a_13623_n4162.n0 a_13623_n4162.n4 1.21355
R16367 a_13623_n4162.n3 a_13623_n4162.n2 0.82773
R16368 a_13623_n4162.n4 a_13623_n4162.n1 0.8005
R16369 a_13623_n4162.n3 a_13623_n4162.n12 0.630329
R16370 a_11023_n9518.n21 a_11023_n9518.t22 56.0276
R16371 a_11023_n9518.n10 a_11023_n9518.t25 56.019
R16372 a_11023_n9518.n12 a_11023_n9518.t30 55.9719
R16373 a_11023_n9518.n6 a_11023_n9518.t20 55.9719
R16374 a_11023_n9518.n14 a_11023_n9518.t35 55.9719
R16375 a_11023_n9518.n5 a_11023_n9518.t27 55.9719
R16376 a_11023_n9518.n16 a_11023_n9518.t36 55.9719
R16377 a_11023_n9518.n4 a_11023_n9518.t32 55.9719
R16378 a_11023_n9518.n17 a_11023_n9518.t23 55.9719
R16379 a_11023_n9518.n2 a_11023_n9518.t37 55.9719
R16380 a_11023_n9518.n22 a_11023_n9518.t34 55.9719
R16381 a_11023_n9518.n10 a_11023_n9518.t31 55.9719
R16382 a_11023_n9518.n10 a_11023_n9518.t39 55.9719
R16383 a_11023_n9518.n9 a_11023_n9518.t26 55.9719
R16384 a_11023_n9518.n9 a_11023_n9518.t33 55.9719
R16385 a_11023_n9518.n7 a_11023_n9518.t21 55.9719
R16386 a_11023_n9518.n7 a_11023_n9518.t28 55.9719
R16387 a_11023_n9518.n8 a_11023_n9518.t24 55.9719
R16388 a_11023_n9518.n8 a_11023_n9518.t29 55.9719
R16389 a_11023_n9518.n27 a_11023_n9518.t38 55.9719
R16390 a_11023_n9518.n12 a_11023_n9518.n11 0.0590857
R16391 a_11023_n9518.n24 a_11023_n9518.n23 4.5005
R16392 a_11023_n9518.n25 a_11023_n9518.n2 4.5005
R16393 a_11023_n9518.n17 a_11023_n9518.n26 4.5005
R16394 a_11023_n9518.n3 a_11023_n9518.n0 4.5005
R16395 a_11023_n9518.n1 a_11023_n9518.n4 4.5005
R16396 a_11023_n9518.n16 a_11023_n9518.n15 4.5005
R16397 a_11023_n9518.n33 a_11023_n9518.n32 4.5005
R16398 a_11023_n9518.n31 a_11023_n9518.n5 4.5005
R16399 a_11023_n9518.n14 a_11023_n9518.n13 4.5005
R16400 a_11023_n9518.n30 a_11023_n9518.n29 4.5005
R16401 a_11023_n9518.n28 a_11023_n9518.n6 4.5005
R16402 a_11023_n9518.n39 a_11023_n9518.n38 3.87048
R16403 a_11023_n9518.n39 a_11023_n9518.n37 3.68704
R16404 a_11023_n9518.n40 a_11023_n9518.n36 3.68704
R16405 a_11023_n9518.n41 a_11023_n9518.n35 3.68704
R16406 a_11023_n9518.n42 a_11023_n9518.n34 3.68704
R16407 a_11023_n9518.n20 a_11023_n9518.n18 3.53719
R16408 a_11023_n9518.n45 a_11023_n9518.n44 3.37808
R16409 a_11023_n9518.n47 a_11023_n9518.n46 3.37808
R16410 a_11023_n9518.n20 a_11023_n9518.n19 3.37808
R16411 a_11023_n9518.n49 a_11023_n9518.n48 3.37783
R16412 a_11023_n9518.n43 a_11023_n9518.n1 1.89107
R16413 a_11023_n9518.n24 a_11023_n9518.n21 1.15666
R16414 a_11023_n9518.n44 a_11023_n9518.t13 0.6505
R16415 a_11023_n9518.n44 a_11023_n9518.t11 0.6505
R16416 a_11023_n9518.n46 a_11023_n9518.t10 0.6505
R16417 a_11023_n9518.n46 a_11023_n9518.t17 0.6505
R16418 a_11023_n9518.n19 a_11023_n9518.t16 0.6505
R16419 a_11023_n9518.n19 a_11023_n9518.t12 0.6505
R16420 a_11023_n9518.n18 a_11023_n9518.t14 0.6505
R16421 a_11023_n9518.n18 a_11023_n9518.t18 0.6505
R16422 a_11023_n9518.t19 a_11023_n9518.n49 0.6505
R16423 a_11023_n9518.n49 a_11023_n9518.t15 0.6505
R16424 a_11023_n9518.n38 a_11023_n9518.t9 0.5855
R16425 a_11023_n9518.n38 a_11023_n9518.t3 0.5855
R16426 a_11023_n9518.n37 a_11023_n9518.t7 0.5855
R16427 a_11023_n9518.n37 a_11023_n9518.t0 0.5855
R16428 a_11023_n9518.n36 a_11023_n9518.t4 0.5855
R16429 a_11023_n9518.n36 a_11023_n9518.t1 0.5855
R16430 a_11023_n9518.n35 a_11023_n9518.t5 0.5855
R16431 a_11023_n9518.n35 a_11023_n9518.t8 0.5855
R16432 a_11023_n9518.n34 a_11023_n9518.t2 0.5855
R16433 a_11023_n9518.n34 a_11023_n9518.t6 0.5855
R16434 a_11023_n9518.n43 a_11023_n9518.n42 0.41138
R16435 a_11023_n9518.n45 a_11023_n9518.n43 0.373278
R16436 a_11023_n9518.n40 a_11023_n9518.n39 0.183939
R16437 a_11023_n9518.n41 a_11023_n9518.n40 0.183939
R16438 a_11023_n9518.n42 a_11023_n9518.n41 0.183939
R16439 a_11023_n9518.n48 a_11023_n9518.n20 0.159616
R16440 a_11023_n9518.n48 a_11023_n9518.n47 0.159616
R16441 a_11023_n9518.n47 a_11023_n9518.n45 0.159616
R16442 a_11023_n9518.n22 a_11023_n9518.n21 0.121859
R16443 a_11023_n9518.n23 a_11023_n9518.n22 0.11975
R16444 a_11023_n9518.n17 a_11023_n9518.n2 0.11975
R16445 a_11023_n9518.n4 a_11023_n9518.n16 0.11975
R16446 a_11023_n9518.n5 a_11023_n9518.n14 0.11975
R16447 a_11023_n9518.n6 a_11023_n9518.n12 0.11975
R16448 a_11023_n9518.n25 a_11023_n9518.n24 0.11975
R16449 a_11023_n9518.n26 a_11023_n9518.n25 0.11975
R16450 a_11023_n9518.n26 a_11023_n9518.n0 0.11975
R16451 a_11023_n9518.n1 a_11023_n9518.n15 0.11975
R16452 a_11023_n9518.n32 a_11023_n9518.n15 0.11975
R16453 a_11023_n9518.n32 a_11023_n9518.n31 0.11975
R16454 a_11023_n9518.n31 a_11023_n9518.n13 0.11975
R16455 a_11023_n9518.n29 a_11023_n9518.n13 0.11975
R16456 a_11023_n9518.n29 a_11023_n9518.n28 0.11975
R16457 a_11023_n9518.n28 a_11023_n9518.n11 2.37025
R16458 a_11023_n9518.n3 a_11023_n9518.n17 0.11975
R16459 a_11023_n9518.n16 a_11023_n9518.n33 0.11975
R16460 a_11023_n9518.n14 a_11023_n9518.n30 0.11975
R16461 a_11023_n9518.n11 a_11023_n9518.n27 1.35571
R16462 a_11023_n9518.n30 a_11023_n9518.n6 0.11975
R16463 a_11023_n9518.n33 a_11023_n9518.n5 0.11975
R16464 a_11023_n9518.n4 a_11023_n9518.n3 0.11975
R16465 a_11023_n9518.n23 a_11023_n9518.n2 0.11975
R16466 a_11023_n9518.n1 a_11023_n9518.n0 0.11975
R16467 a_11023_n9518.n9 a_11023_n9518.n10 0.0946176
R16468 a_11023_n9518.n7 a_11023_n9518.n9 0.0946176
R16469 a_11023_n9518.n8 a_11023_n9518.n7 0.0946176
R16470 a_11023_n9518.n27 a_11023_n9518.n8 0.0946176
R16471 a_23072_n13432.t83 a_23072_n13432.t63 254.709
R16472 a_23072_n13432.t13 a_23072_n13432.t58 254.709
R16473 a_23072_n13432.t37 a_23072_n13432.t97 254.709
R16474 a_23072_n13432.t84 a_23072_n13432.t65 254.709
R16475 a_23072_n13432.t91 a_23072_n13432.t103 254.709
R16476 a_23072_n13432.t10 a_23072_n13432.t93 254.709
R16477 a_23072_n13432.t38 a_23072_n13432.t98 254.709
R16478 a_23072_n13432.t85 a_23072_n13432.t23 254.709
R16479 a_23072_n13432.t30 a_23072_n13432.t94 254.709
R16480 a_23072_n13432.t49 a_23072_n13432.t9 254.709
R16481 a_23072_n13432.t11 a_23072_n13432.t75 254.709
R16482 a_23072_n13432.t67 a_23072_n13432.t39 254.709
R16483 a_23072_n13432.t59 a_23072_n13432.t79 254.709
R16484 a_23072_n13432.t68 a_23072_n13432.t21 254.709
R16485 a_23072_n13432.t45 a_23072_n13432.t66 254.709
R16486 a_23072_n13432.t101 a_23072_n13432.t53 196.517
R16487 a_23072_n13432.n50 a_23072_n13432.t81 31.4493
R16488 a_23072_n13432.n44 a_23072_n13432.t34 31.4493
R16489 a_23072_n13432.n39 a_23072_n13432.t62 31.4493
R16490 a_23072_n13432.n36 a_23072_n13432.t14 31.4493
R16491 a_23072_n13432.n33 a_23072_n13432.t69 31.4493
R16492 a_23072_n13432.n29 a_23072_n13432.t57 31.4493
R16493 a_23072_n13432.n37 a_23072_n13432.t73 31.4493
R16494 a_23072_n13432.n25 a_23072_n13432.t77 31.4493
R16495 a_23072_n13432.n26 a_23072_n13432.t48 31.4493
R16496 a_23072_n13432.n43 a_23072_n13432.t50 31.4493
R16497 a_23072_n13432.n45 a_23072_n13432.t19 31.4493
R16498 a_23072_n13432.n47 a_23072_n13432.t41 31.4493
R16499 a_23072_n13432.n19 a_23072_n13432.t35 31.4493
R16500 a_23072_n13432.n18 a_23072_n13432.t61 31.4493
R16501 a_23072_n13432.n17 a_23072_n13432.t102 31.4493
R16502 a_23072_n13432.n27 a_23072_n13432.n25 29.66
R16503 a_23072_n13432.t63 a_23072_n13432.t36 23.7012
R16504 a_23072_n13432.t58 a_23072_n13432.t12 23.7012
R16505 a_23072_n13432.t97 a_23072_n13432.t24 23.7012
R16506 a_23072_n13432.t65 a_23072_n13432.t82 23.7012
R16507 a_23072_n13432.t103 a_23072_n13432.t18 23.7012
R16508 a_23072_n13432.t93 a_23072_n13432.t95 23.7012
R16509 a_23072_n13432.t98 a_23072_n13432.t25 23.7012
R16510 a_23072_n13432.t23 a_23072_n13432.t29 23.7012
R16511 a_23072_n13432.t94 a_23072_n13432.t26 23.7012
R16512 a_23072_n13432.t9 a_23072_n13432.t70 23.7012
R16513 a_23072_n13432.t75 a_23072_n13432.t47 23.7012
R16514 a_23072_n13432.t39 a_23072_n13432.t31 23.7012
R16515 a_23072_n13432.t79 a_23072_n13432.t55 23.7012
R16516 a_23072_n13432.t21 a_23072_n13432.t99 23.7012
R16517 a_23072_n13432.t66 a_23072_n13432.t40 23.7012
R16518 a_23072_n13432.t53 a_23072_n13432.t43 23.4396
R16519 a_23072_n13432.n16 a_23072_n13432.n14 22.364
R16520 a_23072_n13432.n2 a_23072_n13432.n17 18.725
R16521 a_23072_n13432.n48 a_23072_n13432.n47 18.005
R16522 a_23072_n13432.n34 a_23072_n13432.n33 17.865
R16523 a_23072_n13432.n6 a_23072_n13432.n43 17.825
R16524 a_23072_n13432.n8 a_23072_n13432.n50 17.285
R16525 a_23072_n13432.n30 a_23072_n13432.n29 17.285
R16526 a_23072_n13432.n0 a_23072_n13432.n21 17.0555
R16527 a_23072_n13432.n1 a_23072_n13432.n16 16.3355
R16528 a_23072_n13432.n30 a_23072_n13432.n28 15.6981
R16529 a_23072_n13432.n35 a_23072_n13432.t86 14.2998
R16530 a_23072_n13432.n35 a_23072_n13432.t101 13.8705
R16531 a_23072_n13432.n46 a_23072_n13432.n45 13.145
R16532 a_23072_n13432.n27 a_23072_n13432.n26 12.965
R16533 a_23072_n13432.n7 a_23072_n13432.n40 12.9155
R16534 a_23072_n13432.n5 a_23072_n13432.n36 12.785
R16535 a_23072_n13432.n38 a_23072_n13432.n37 12.7763
R16536 a_23072_n13432.n5 a_23072_n13432.n35 12.6959
R16537 a_23072_n13432.n7 a_23072_n13432.n44 12.645
R16538 a_23072_n13432.n40 a_23072_n13432.n39 12.645
R16539 a_23072_n13432.n4 a_23072_n13432.n18 12.645
R16540 a_23072_n13432.n11 a_23072_n13432.n19 12.5963
R16541 a_23072_n13432.n22 a_23072_n13432.n20 12.3305
R16542 a_23072_n13432.n6 a_23072_n13432.n42 12.2781
R16543 a_23072_n13432.n4 a_23072_n13432.n2 11.3855
R16544 a_23072_n13432.n2 a_23072_n13432.n13 10.6013
R16545 a_23072_n13432.n6 a_23072_n13432.n41 10.0805
R16546 a_23072_n13432.n12 a_23072_n13432.n24 9.9005
R16547 a_23072_n13432.n22 a_23072_n13432.n0 9.7205
R16548 a_23072_n13432.n1 a_23072_n13432.t76 9.70587
R16549 a_23072_n13432.n12 a_23072_n13432.n38 9.4955
R16550 a_23072_n13432.n2 a_23072_n13432.n1 9.3605
R16551 a_23072_n13432.n32 a_23072_n13432.n31 9.0005
R16552 a_23072_n13432.n8 a_23072_n13432.n11 8.9555
R16553 a_23072_n13432.n4 a_23072_n13432.n8 8.1005
R16554 a_23072_n13432.n48 a_23072_n13432.n46 8.0555
R16555 a_23072_n13432.n5 a_23072_n13432.n34 7.4255
R16556 a_23072_n13432.n4 a_23072_n13432.n3 7.2905
R16557 a_23072_n13432.n9 a_23072_n13432.t2 7.13263
R16558 a_23072_n13432.n9 a_23072_n13432.t3 7.13263
R16559 a_23072_n13432.n49 a_23072_n13432.n23 6.7955
R16560 a_23072_n13432.n50 a_23072_n13432.t83 6.79462
R16561 a_23072_n13432.n44 a_23072_n13432.t13 6.79462
R16562 a_23072_n13432.n39 a_23072_n13432.t37 6.79462
R16563 a_23072_n13432.n36 a_23072_n13432.t84 6.79462
R16564 a_23072_n13432.n33 a_23072_n13432.t91 6.79462
R16565 a_23072_n13432.n29 a_23072_n13432.t10 6.79462
R16566 a_23072_n13432.n37 a_23072_n13432.t38 6.79462
R16567 a_23072_n13432.n25 a_23072_n13432.t85 6.79462
R16568 a_23072_n13432.n26 a_23072_n13432.t30 6.79462
R16569 a_23072_n13432.n43 a_23072_n13432.t49 6.79462
R16570 a_23072_n13432.n45 a_23072_n13432.t11 6.79462
R16571 a_23072_n13432.n47 a_23072_n13432.t67 6.79462
R16572 a_23072_n13432.n19 a_23072_n13432.t59 6.79462
R16573 a_23072_n13432.n18 a_23072_n13432.t68 6.79462
R16574 a_23072_n13432.n17 a_23072_n13432.t45 6.79462
R16575 a_23072_n13432.n32 a_23072_n13432.n30 6.7505
R16576 a_23072_n13432.n41 a_23072_n13432.t46 6.71423
R16577 a_23072_n13432.n23 a_23072_n13432.t56 6.71423
R16578 a_23072_n13432.n10 a_23072_n13432.t74 6.71423
R16579 a_23072_n13432.n3 a_23072_n13432.t8 6.71423
R16580 a_23072_n13432.n1 a_23072_n13432.t80 6.71423
R16581 a_23072_n13432.n14 a_23072_n13432.t64 6.71423
R16582 a_23072_n13432.n24 a_23072_n13432.t52 6.56378
R16583 a_23072_n13432.n0 a_23072_n13432.t16 6.56378
R16584 a_23072_n13432.n21 a_23072_n13432.t89 6.56378
R16585 a_23072_n13432.n49 a_23072_n13432.n48 6.4805
R16586 a_23072_n13432.n9 a_23072_n13432.t4 6.43746
R16587 a_23072_n13432.n9 a_23072_n13432.t1 6.43746
R16588 a_23072_n13432.n9 a_23072_n13432.n4 6.4355
R16589 a_23072_n13432.n31 a_23072_n13432.t42 6.41334
R16590 a_23072_n13432.n20 a_23072_n13432.t92 6.41334
R16591 a_23072_n13432.n51 a_23072_n13432.t78 6.3005
R16592 a_23072_n13432.n28 a_23072_n13432.t60 6.3005
R16593 a_23072_n13432.n42 a_23072_n13432.t88 6.3005
R16594 a_23072_n13432.n15 a_23072_n13432.t33 6.3005
R16595 a_23072_n13432.n13 a_23072_n13432.t72 6.3005
R16596 a_23072_n13432.n8 a_23072_n13432.n49 6.2555
R16597 a_23072_n13432.n40 a_23072_n13432.n12 6.2555
R16598 a_23072_n13432.n12 a_23072_n13432.n27 6.2105
R16599 a_23072_n13432.n11 a_23072_n13432.n10 6.0755
R16600 a_23072_n13432.n38 a_23072_n13432.n5 5.6705
R16601 a_23072_n13432.n51 a_23072_n13432.t90 5.6196
R16602 a_23072_n13432.n28 a_23072_n13432.t71 5.6196
R16603 a_23072_n13432.n42 a_23072_n13432.t96 5.6196
R16604 a_23072_n13432.n15 a_23072_n13432.t28 5.6196
R16605 a_23072_n13432.n13 a_23072_n13432.t44 5.6196
R16606 a_23072_n13432.n34 a_23072_n13432.n32 5.5805
R16607 a_23072_n13432.n31 a_23072_n13432.t87 5.50677
R16608 a_23072_n13432.n20 a_23072_n13432.t20 5.50677
R16609 a_23072_n13432.n9 a_23072_n13432.t7 5.41151
R16610 a_23072_n13432.n24 a_23072_n13432.t54 5.35632
R16611 a_23072_n13432.n0 a_23072_n13432.t51 5.35632
R16612 a_23072_n13432.n21 a_23072_n13432.t22 5.35632
R16613 a_23072_n13432.n7 a_23072_n13432.n6 5.2205
R16614 a_23072_n13432.n41 a_23072_n13432.t32 5.20587
R16615 a_23072_n13432.n23 a_23072_n13432.t15 5.20587
R16616 a_23072_n13432.n10 a_23072_n13432.t100 5.20587
R16617 a_23072_n13432.n3 a_23072_n13432.t17 5.20587
R16618 a_23072_n13432.n14 a_23072_n13432.t27 5.20587
R16619 a_23072_n13432.n9 a_23072_n13432.t6 4.86588
R16620 a_23072_n13432.n9 a_23072_n13432.t5 4.78151
R16621 a_23072_n13432.n46 a_23072_n13432.n7 4.7255
R16622 a_23072_n13432.n11 a_23072_n13432.n22 4.6805
R16623 a_23072_n13432.t0 a_23072_n13432.n9 4.63548
R16624 a_23072_n13432.n4 a_23072_n13432.n51 4.53811
R16625 a_23072_n13432.n16 a_23072_n13432.n15 4.53811
R16626 a_29920_n3900.n12 a_29920_n3900.n9 38.8088
R16627 a_29920_n3900.n5 a_29920_n3900.t13 29.2005
R16628 a_29920_n3900.n13 a_29920_n3900.t22 23.0685
R16629 a_29920_n3900.n0 a_29920_n3900.n5 21.5736
R16630 a_29920_n3900.n9 a_29920_n3900.t21 18.9805
R16631 a_29920_n3900.n14 a_29920_n3900.t4 17.2042
R16632 a_29920_n3900.n14 a_29920_n3900.t6 16.6445
R16633 a_29920_n3900.n1 a_29920_n3900.n2 4.45624
R16634 a_29920_n3900.n11 a_29920_n3900.t11 16.4255
R16635 a_29920_n3900.n1 a_29920_n3900.t12 16.4255
R16636 a_29920_n3900.n10 a_29920_n3900.t20 16.4255
R16637 a_29920_n3900.n4 a_29920_n3900.t15 16.4012
R16638 a_29920_n3900.n11 a_29920_n3900.t3 16.3282
R16639 a_29920_n3900.n10 a_29920_n3900.t9 16.3282
R16640 a_29920_n3900.n7 a_29920_n3900.t14 15.8415
R16641 a_29920_n3900.n6 a_29920_n3900.t17 15.8415
R16642 a_29920_n3900.n8 a_29920_n3900.t10 15.8415
R16643 a_29920_n3900.n1 a_29920_n3900.t5 14.7952
R16644 a_29920_n3900.n0 a_29920_n3900.n8 13.5501
R16645 a_29920_n3900.n4 a_29920_n3900.t8 13.4447
R16646 a_29920_n3900.n5 a_29920_n3900.t18 12.1428
R16647 a_29920_n3900.n9 a_29920_n3900.t16 11.4372
R16648 a_29920_n3900.n7 a_29920_n3900.t7 11.3763
R16649 a_29920_n3900.n6 a_29920_n3900.t2 11.3763
R16650 a_29920_n3900.n8 a_29920_n3900.t23 11.3763
R16651 a_29920_n3900.n16 a_29920_n3900.n12 10.9805
R16652 a_29920_n3900.n13 a_29920_n3900.t19 10.7802
R16653 a_29920_n3900.n8 a_29920_n3900.n6 10.5449
R16654 a_29920_n3900.n8 a_29920_n3900.n7 10.5449
R16655 a_29920_n3900.n3 a_29920_n3900.n2 2.5054
R16656 a_29920_n3900.n4 a_29920_n3900.n2 4.33683
R16657 a_29920_n3900.n17 a_29920_n3900.n0 9.0005
R16658 a_29920_n3900.n0 a_29920_n3900.n16 8.8205
R16659 a_29920_n3900.n3 a_29920_n3900.n10 8.79675
R16660 a_29920_n3900.n15 a_29920_n3900.n14 8.64897
R16661 a_29920_n3900.n15 a_29920_n3900.n13 8.33894
R16662 a_29920_n3900.n3 a_29920_n3900.n11 8.04925
R16663 a_29920_n3900.n17 a_29920_n3900.t0 6.6642
R16664 a_29920_n3900.n12 a_29920_n3900.n3 5.5155
R16665 a_29920_n3900.n16 a_29920_n3900.n15 4.5005
R16666 a_29920_n3900.t1 a_29920_n3900.n17 2.88679
R16667 a_21772_n3588.n2 a_21772_n3588.t13 15.8415
R16668 a_21772_n3588.n3 a_21772_n3588.t19 15.8415
R16669 a_21772_n3588.n4 a_21772_n3588.t16 15.8415
R16670 a_21772_n3588.n5 a_21772_n3588.t4 15.8415
R16671 a_21772_n3588.n6 a_21772_n3588.t6 15.8415
R16672 a_21772_n3588.n7 a_21772_n3588.t10 15.8415
R16673 a_21772_n3588.n1 a_21772_n3588.t9 15.8415
R16674 a_21772_n3588.n0 a_21772_n3588.t11 15.8415
R16675 a_21772_n3588.n2 a_21772_n3588.t12 13.4447
R16676 a_21772_n3588.n3 a_21772_n3588.t14 13.4447
R16677 a_21772_n3588.n4 a_21772_n3588.t15 13.4447
R16678 a_21772_n3588.n5 a_21772_n3588.t17 13.4447
R16679 a_21772_n3588.n6 a_21772_n3588.t5 13.4447
R16680 a_21772_n3588.n7 a_21772_n3588.t18 13.4447
R16681 a_21772_n3588.n1 a_21772_n3588.t7 13.4447
R16682 a_21772_n3588.n0 a_21772_n3588.t8 13.4447
R16683 a_21772_n3588.n3 a_21772_n3588.n2 10.5449
R16684 a_21772_n3588.n4 a_21772_n3588.n3 10.5449
R16685 a_21772_n3588.n5 a_21772_n3588.n4 10.5449
R16686 a_21772_n3588.n6 a_21772_n3588.n5 10.5449
R16687 a_21772_n3588.n7 a_21772_n3588.n6 10.5449
R16688 a_21772_n3588.n0 a_21772_n3588.n1 10.5449
R16689 a_21772_n3588.n0 a_21772_n3588.n7 10.5449
R16690 a_21772_n3588.n0 a_21772_n3588.t2 7.22489
R16691 a_21772_n3588.t1 a_21772_n3588.n0 7.12153
R16692 a_21772_n3588.n0 a_21772_n3588.t0 6.36702
R16693 a_21772_n3588.n0 a_21772_n3588.t3 5.62673
R16694 a_13623_n20230.n1 a_13623_n20230.t33 56.1018
R16695 a_13623_n20230.n2 a_13623_n20230.t42 56.0719
R16696 a_13623_n20230.n1 a_13623_n20230.t37 56.0141
R16697 a_13623_n20230.n1 a_13623_n20230.t44 55.9719
R16698 a_13623_n20230.n1 a_13623_n20230.t27 55.9719
R16699 a_13623_n20230.n1 a_13623_n20230.t35 55.9719
R16700 a_13623_n20230.n1 a_13623_n20230.t19 55.9719
R16701 a_13623_n20230.n1 a_13623_n20230.t40 55.9719
R16702 a_13623_n20230.n1 a_13623_n20230.t21 55.9719
R16703 a_13623_n20230.n1 a_13623_n20230.t32 55.9719
R16704 a_13623_n20230.n1 a_13623_n20230.t43 55.9719
R16705 a_13623_n20230.n1 a_13623_n20230.t26 55.9719
R16706 a_13623_n20230.n1 a_13623_n20230.t17 55.9719
R16707 a_13623_n20230.n1 a_13623_n20230.t30 55.9719
R16708 a_13623_n20230.n1 a_13623_n20230.t38 55.9719
R16709 a_13623_n20230.n1 a_13623_n20230.t23 55.9719
R16710 a_13623_n20230.n1 a_13623_n20230.t45 55.9719
R16711 a_13623_n20230.n1 a_13623_n20230.t24 55.9719
R16712 a_13623_n20230.n1 a_13623_n20230.t36 55.9719
R16713 a_13623_n20230.n1 a_13623_n20230.t16 55.9719
R16714 a_13623_n20230.n1 a_13623_n20230.t29 55.9719
R16715 a_13623_n20230.n2 a_13623_n20230.t25 55.9719
R16716 a_13623_n20230.n2 a_13623_n20230.t34 55.9719
R16717 a_13623_n20230.n2 a_13623_n20230.t28 55.9719
R16718 a_13623_n20230.n2 a_13623_n20230.t39 55.9719
R16719 a_13623_n20230.n2 a_13623_n20230.t20 55.9719
R16720 a_13623_n20230.n2 a_13623_n20230.t31 55.9719
R16721 a_13623_n20230.n4 a_13623_n20230.t41 55.9719
R16722 a_13623_n20230.n4 a_13623_n20230.t22 55.9719
R16723 a_13623_n20230.n4 a_13623_n20230.t18 55.9719
R16724 a_13623_n20230.n0 a_13623_n20230.n1 38.7327
R16725 a_13623_n20230.n0 a_13623_n20230.n8 6.90733
R16726 a_13623_n20230.n3 a_13623_n20230.n10 6.89497
R16727 a_13623_n20230.n3 a_13623_n20230.n9 6.3768
R16728 a_13623_n20230.n0 a_13623_n20230.n7 6.3768
R16729 a_13623_n20230.n0 a_13623_n20230.n6 3.21104
R16730 a_13623_n20230.n0 a_13623_n20230.n5 2.7042
R16731 a_13623_n20230.n0 a_13623_n20230.n11 2.7042
R16732 a_13623_n20230.n12 a_13623_n20230.n0 2.7042
R16733 a_13623_n20230.n6 a_13623_n20230.t13 2.06607
R16734 a_13623_n20230.n5 a_13623_n20230.t14 2.06607
R16735 a_13623_n20230.n11 a_13623_n20230.t10 2.06607
R16736 a_13623_n20230.n12 a_13623_n20230.t9 2.06607
R16737 a_13623_n20230.n9 a_13623_n20230.t0 1.99806
R16738 a_13623_n20230.n9 a_13623_n20230.t7 1.99806
R16739 a_13623_n20230.n10 a_13623_n20230.t6 1.99806
R16740 a_13623_n20230.n10 a_13623_n20230.t5 1.99806
R16741 a_13623_n20230.n8 a_13623_n20230.t3 1.99806
R16742 a_13623_n20230.n8 a_13623_n20230.t4 1.99806
R16743 a_13623_n20230.n7 a_13623_n20230.t1 1.99806
R16744 a_13623_n20230.n7 a_13623_n20230.t2 1.99806
R16745 a_13623_n20230.n6 a_13623_n20230.t11 1.4923
R16746 a_13623_n20230.n5 a_13623_n20230.t12 1.4923
R16747 a_13623_n20230.n11 a_13623_n20230.t8 1.4923
R16748 a_13623_n20230.t15 a_13623_n20230.n12 1.4923
R16749 a_13623_n20230.n0 a_13623_n20230.n3 1.35826
R16750 a_13623_n20230.n1 a_13623_n20230.n4 1.21355
R16751 a_13623_n20230.n4 a_13623_n20230.n2 0.8005
R16752 a_25020_n8200.n0 a_25020_n8200.n1 30.5016
R16753 a_25020_n8200.n1 a_25020_n8200.t6 29.2005
R16754 a_25020_n8200.n0 a_25020_n8200.n3 28.2928
R16755 a_25020_n8200.n3 a_25020_n8200.t5 20.1607
R16756 a_25020_n8200.n0 a_25020_n8200.n2 18.2882
R16757 a_25020_n8200.n2 a_25020_n8200.t7 17.5205
R16758 a_25020_n8200.n1 a_25020_n8200.t4 12.1428
R16759 a_25020_n8200.n2 a_25020_n8200.t3 11.5588
R16760 a_25020_n8200.t1 a_25020_n8200.n0 11.5205
R16761 a_25020_n8200.n3 a_25020_n8200.t2 10.8288
R16762 a_25020_n8200.t1 a_25020_n8200.t0 8.55859
R16763 a_4001_4292.n3 a_4001_4292.t6 67.9167
R16764 a_4001_4292.n3 a_4001_4292.t14 65.1645
R16765 a_4001_4292.n0 a_4001_4292.t4 56.1589
R16766 a_4001_4292.n2 a_4001_4292.t12 55.9719
R16767 a_4001_4292.n2 a_4001_4292.t11 55.9719
R16768 a_4001_4292.n1 a_4001_4292.t13 55.9719
R16769 a_4001_4292.n1 a_4001_4292.t10 55.9719
R16770 a_4001_4292.n1 a_4001_4292.t9 55.9719
R16771 a_4001_4292.n1 a_4001_4292.t8 55.9719
R16772 a_4001_4292.n0 a_4001_4292.t7 55.9719
R16773 a_4001_4292.n0 a_4001_4292.t3 55.9719
R16774 a_4001_4292.n0 a_4001_4292.t5 55.9719
R16775 a_4001_4292.n3 a_4001_4292.n2 13.3524
R16776 a_4001_4292.n4 a_4001_4292.n3 9.7565
R16777 a_4001_4292.n5 a_4001_4292.t2 3.69547
R16778 a_4001_4292.t1 a_4001_4292.n5 3.12815
R16779 a_4001_4292.n4 a_4001_4292.t0 2.88322
R16780 a_4001_4292.n5 a_4001_4292.n4 1.535
R16781 a_4001_4292.n1 a_4001_4292.n0 0.748552
R16782 a_4001_4292.n2 a_4001_4292.n1 0.748552
R16783 a_13501_n14494.n1 a_13501_n14494.t2 15.8618
R16784 a_13501_n14494.n0 a_13501_n14494.t3 15.8393
R16785 a_13501_n14494.n1 a_13501_n14494.t16 15.7537
R16786 a_13501_n14494.n0 a_13501_n14494.t15 15.7496
R16787 a_13501_n14494.n0 a_13501_n14494.n2 14.963
R16788 a_13501_n14494.n1 a_13501_n14494.n4 14.9583
R16789 a_13501_n14494.n1 a_13501_n14494.n7 14.9559
R16790 a_13501_n14494.n1 a_13501_n14494.n8 14.9547
R16791 a_13501_n14494.n0 a_13501_n14494.n3 14.7096
R16792 a_13501_n14494.n9 a_13501_n14494.n1 14.7035
R16793 a_13501_n14494.n1 a_13501_n14494.n5 14.7035
R16794 a_13501_n14494.n1 a_13501_n14494.n6 14.6941
R16795 a_13501_n14494.n6 a_13501_n14494.t19 0.6505
R16796 a_13501_n14494.n6 a_13501_n14494.t12 0.6505
R16797 a_13501_n14494.n5 a_13501_n14494.t10 0.6505
R16798 a_13501_n14494.n5 a_13501_n14494.t14 0.6505
R16799 a_13501_n14494.n3 a_13501_n14494.t13 0.6505
R16800 a_13501_n14494.n3 a_13501_n14494.t17 0.6505
R16801 a_13501_n14494.t18 a_13501_n14494.n9 0.6505
R16802 a_13501_n14494.n9 a_13501_n14494.t11 0.6505
R16803 a_13501_n14494.n7 a_13501_n14494.t9 0.5855
R16804 a_13501_n14494.n7 a_13501_n14494.t6 0.5855
R16805 a_13501_n14494.n8 a_13501_n14494.t0 0.5855
R16806 a_13501_n14494.n8 a_13501_n14494.t7 0.5855
R16807 a_13501_n14494.n4 a_13501_n14494.t8 0.5855
R16808 a_13501_n14494.n4 a_13501_n14494.t4 0.5855
R16809 a_13501_n14494.n2 a_13501_n14494.t5 0.5855
R16810 a_13501_n14494.n2 a_13501_n14494.t1 0.5855
R16811 a_13501_n14494.n1 a_13501_n14494.n0 0.158862
R16812 a_33776_n5896.n9 a_33776_n5896.t20 15.7685
R16813 a_33776_n5896.n10 a_33776_n5896.t11 15.7685
R16814 a_33776_n5896.n3 a_33776_n5896.t17 15.7685
R16815 a_33776_n5896.n4 a_33776_n5896.t9 15.7685
R16816 a_33776_n5896.n5 a_33776_n5896.t19 15.7685
R16817 a_33776_n5896.n6 a_33776_n5896.t8 15.7685
R16818 a_33776_n5896.n7 a_33776_n5896.t15 15.7685
R16819 a_33776_n5896.n8 a_33776_n5896.t18 15.7685
R16820 a_33776_n5896.n9 a_33776_n5896.t10 11.6197
R16821 a_33776_n5896.n10 a_33776_n5896.t22 11.6197
R16822 a_33776_n5896.n3 a_33776_n5896.t14 11.6197
R16823 a_33776_n5896.n4 a_33776_n5896.t13 11.6197
R16824 a_33776_n5896.n5 a_33776_n5896.t16 11.6197
R16825 a_33776_n5896.n6 a_33776_n5896.t12 11.6197
R16826 a_33776_n5896.n7 a_33776_n5896.t21 11.6197
R16827 a_33776_n5896.n8 a_33776_n5896.t7 11.6197
R16828 a_33776_n5896.n10 a_33776_n5896.n9 10.5449
R16829 a_33776_n5896.n4 a_33776_n5896.n3 10.5449
R16830 a_33776_n5896.n5 a_33776_n5896.n4 10.5449
R16831 a_33776_n5896.n6 a_33776_n5896.n5 10.5449
R16832 a_33776_n5896.n7 a_33776_n5896.n6 10.5449
R16833 a_33776_n5896.n8 a_33776_n5896.n7 10.5449
R16834 a_33776_n5896.n0 a_33776_n5896.t0 10.4819
R16835 a_33776_n5896.n11 a_33776_n5896.n8 8.41578
R16836 a_33776_n5896.n0 a_33776_n5896.n2 7.31398
R16837 a_33776_n5896.n12 a_33776_n5896.n0 6.25311
R16838 a_33776_n5896.n0 a_33776_n5896.n1 5.37659
R16839 a_33776_n5896.n2 a_33776_n5896.t1 4.04494
R16840 a_33776_n5896.n2 a_33776_n5896.t2 4.04494
R16841 a_33776_n5896.n1 a_33776_n5896.t5 3.07367
R16842 a_33776_n5896.n1 a_33776_n5896.t3 3.07367
R16843 a_33776_n5896.t6 a_33776_n5896.n12 3.07367
R16844 a_33776_n5896.n12 a_33776_n5896.t4 3.07367
R16845 a_33776_n5896.n0 a_33776_n5896.n11 2.93567
R16846 a_33776_n5896.n11 a_33776_n5896.n10 2.12967
R16847 a_34708_n5896.n10 a_34708_n5896.t27 31.6987
R16848 a_34708_n5896.n16 a_34708_n5896.t17 31.6987
R16849 a_34708_n5896.n11 a_34708_n5896.t29 18.6885
R16850 a_34708_n5896.n12 a_34708_n5896.t25 18.6885
R16851 a_34708_n5896.n10 a_34708_n5896.t20 18.6885
R16852 a_34708_n5896.n16 a_34708_n5896.t28 18.6885
R16853 a_34708_n5896.n14 a_34708_n5896.t16 18.6885
R16854 a_34708_n5896.n15 a_34708_n5896.t19 18.6885
R16855 a_34708_n5896.n11 a_34708_n5896.t21 11.1938
R16856 a_34708_n5896.n12 a_34708_n5896.t18 11.1938
R16857 a_34708_n5896.n10 a_34708_n5896.t26 11.1938
R16858 a_34708_n5896.n16 a_34708_n5896.t23 11.1938
R16859 a_34708_n5896.n14 a_34708_n5896.t24 11.1938
R16860 a_34708_n5896.n15 a_34708_n5896.t22 11.1938
R16861 a_34708_n5896.n12 a_34708_n5896.n11 10.5449
R16862 a_34708_n5896.n15 a_34708_n5896.n14 10.5449
R16863 a_34708_n5896.n18 a_34708_n5896.n17 9.36336
R16864 a_34708_n5896.n18 a_34708_n5896.n13 7.21225
R16865 a_34708_n5896.n0 a_34708_n5896.n9 7.13263
R16866 a_34708_n5896.n2 a_34708_n5896.n7 7.13263
R16867 a_34708_n5896.n13 a_34708_n5896.n10 6.48939
R16868 a_34708_n5896.n17 a_34708_n5896.n16 6.48939
R16869 a_34708_n5896.n0 a_34708_n5896.n8 6.43746
R16870 a_34708_n5896.n2 a_34708_n5896.n6 6.43746
R16871 a_34708_n5896.n1 a_34708_n5896.n18 4.5005
R16872 a_34708_n5896.n13 a_34708_n5896.n12 4.05606
R16873 a_34708_n5896.n17 a_34708_n5896.n15 4.05606
R16874 a_34708_n5896.n9 a_34708_n5896.t3 3.8098
R16875 a_34708_n5896.n9 a_34708_n5896.t4 3.8098
R16876 a_34708_n5896.n8 a_34708_n5896.t2 3.8098
R16877 a_34708_n5896.n8 a_34708_n5896.t5 3.8098
R16878 a_34708_n5896.n6 a_34708_n5896.t1 3.8098
R16879 a_34708_n5896.n6 a_34708_n5896.t7 3.8098
R16880 a_34708_n5896.n7 a_34708_n5896.t0 3.8098
R16881 a_34708_n5896.n7 a_34708_n5896.t6 3.8098
R16882 a_34708_n5896.n1 a_34708_n5896.n5 3.34593
R16883 a_34708_n5896.n1 a_34708_n5896.n3 3.34593
R16884 a_34708_n5896.n1 a_34708_n5896.n4 2.71593
R16885 a_34708_n5896.n19 a_34708_n5896.n1 2.71593
R16886 a_34708_n5896.n5 a_34708_n5896.t13 2.06607
R16887 a_34708_n5896.n5 a_34708_n5896.t8 2.06607
R16888 a_34708_n5896.n4 a_34708_n5896.t12 2.06607
R16889 a_34708_n5896.n4 a_34708_n5896.t10 2.06607
R16890 a_34708_n5896.n3 a_34708_n5896.t11 2.06607
R16891 a_34708_n5896.n3 a_34708_n5896.t14 2.06607
R16892 a_34708_n5896.n19 a_34708_n5896.t9 2.06607
R16893 a_34708_n5896.t15 a_34708_n5896.n19 2.06607
R16894 a_34708_n5896.n1 a_34708_n5896.n0 0.797178
R16895 a_34708_n5896.n0 a_34708_n5896.n2 0.577741
R16896 a_29076_n8292.n5 a_29076_n8292.n4 25.2911
R16897 a_29076_n8292.n7 a_29076_n8292.n6 21.8536
R16898 a_29076_n8292.n2 a_29076_n8292.t4 19.5645
R16899 a_29076_n8292.n6 a_29076_n8292.t11 19.5523
R16900 a_29076_n8292.n2 a_29076_n8292.t10 18.4938
R16901 a_29076_n8292.n4 a_29076_n8292.t6 17.4475
R16902 a_29076_n8292.n1 a_29076_n8292.t7 16.7662
R16903 a_29076_n8292.n1 a_29076_n8292.t9 14.3815
R16904 a_29076_n8292.n4 a_29076_n8292.t8 12.7755
R16905 a_29076_n8292.n7 a_29076_n8292.n5 11.0705
R16906 a_29076_n8292.n0 a_29076_n8292.n7 10.6205
R16907 a_29076_n8292.n6 a_29076_n8292.t5 9.79467
R16908 a_29076_n8292.n3 a_29076_n8292.n2 9.20964
R16909 a_29076_n8292.n5 a_29076_n8292.n3 8.9105
R16910 a_29076_n8292.n3 a_29076_n8292.n1 8.15261
R16911 a_29076_n8292.n0 a_29076_n8292.t2 7.76131
R16912 a_29076_n8292.t1 a_29076_n8292.n0 6.44627
R16913 a_29076_n8292.n0 a_29076_n8292.t0 5.98178
R16914 a_29076_n8292.n0 a_29076_n8292.t3 5.2005
R16915 a_21996_332.n0 a_21996_332.n1 59.4642
R16916 a_21996_332.n1 a_21996_332.t2 18.141
R16917 a_21996_332.n1 a_21996_332.t3 11.863
R16918 a_21996_332.n0 a_21996_332.t0 8.56922
R16919 a_21996_332.t1 a_21996_332.n0 4.8813
R16920 a_13501_n17172.n1 a_13501_n17172.t0 15.8618
R16921 a_13501_n17172.n0 a_13501_n17172.t9 15.8393
R16922 a_13501_n17172.t18 a_13501_n17172.n1 15.7537
R16923 a_13501_n17172.n0 a_13501_n17172.t17 15.7496
R16924 a_13501_n17172.n0 a_13501_n17172.n2 14.963
R16925 a_13501_n17172.n1 a_13501_n17172.n4 14.9583
R16926 a_13501_n17172.n1 a_13501_n17172.n8 14.9559
R16927 a_13501_n17172.n1 a_13501_n17172.n7 14.9547
R16928 a_13501_n17172.n0 a_13501_n17172.n3 14.7096
R16929 a_13501_n17172.n1 a_13501_n17172.n6 14.7035
R16930 a_13501_n17172.n1 a_13501_n17172.n5 14.7035
R16931 a_13501_n17172.n1 a_13501_n17172.n9 14.6941
R16932 a_13501_n17172.n9 a_13501_n17172.t11 0.6505
R16933 a_13501_n17172.n9 a_13501_n17172.t14 0.6505
R16934 a_13501_n17172.n6 a_13501_n17172.t10 0.6505
R16935 a_13501_n17172.n6 a_13501_n17172.t13 0.6505
R16936 a_13501_n17172.n5 a_13501_n17172.t12 0.6505
R16937 a_13501_n17172.n5 a_13501_n17172.t16 0.6505
R16938 a_13501_n17172.n3 a_13501_n17172.t15 0.6505
R16939 a_13501_n17172.n3 a_13501_n17172.t19 0.6505
R16940 a_13501_n17172.n8 a_13501_n17172.t3 0.5855
R16941 a_13501_n17172.n8 a_13501_n17172.t6 0.5855
R16942 a_13501_n17172.n7 a_13501_n17172.t2 0.5855
R16943 a_13501_n17172.n7 a_13501_n17172.t5 0.5855
R16944 a_13501_n17172.n4 a_13501_n17172.t4 0.5855
R16945 a_13501_n17172.n4 a_13501_n17172.t8 0.5855
R16946 a_13501_n17172.n2 a_13501_n17172.t7 0.5855
R16947 a_13501_n17172.n2 a_13501_n17172.t1 0.5855
R16948 a_13501_n17172.n1 a_13501_n17172.n0 0.158862
R16949 a_3935_4156.n3 a_3935_4156.t9 68.0895
R16950 a_3935_4156.n3 a_3935_4156.t8 65.1645
R16951 a_3935_4156.n0 a_3935_4156.t13 56.1655
R16952 a_3935_4156.n2 a_3935_4156.t3 55.9719
R16953 a_3935_4156.n2 a_3935_4156.t12 55.9719
R16954 a_3935_4156.n1 a_3935_4156.t10 55.9719
R16955 a_3935_4156.n1 a_3935_4156.t6 55.9719
R16956 a_3935_4156.n1 a_3935_4156.t11 55.9719
R16957 a_3935_4156.n1 a_3935_4156.t7 55.9719
R16958 a_3935_4156.n0 a_3935_4156.t5 55.9719
R16959 a_3935_4156.n0 a_3935_4156.t4 55.9719
R16960 a_3935_4156.n0 a_3935_4156.t14 55.9719
R16961 a_3935_4156.n3 a_3935_4156.n2 26.3688
R16962 a_3935_4156.n4 a_3935_4156.n3 9.8735
R16963 a_3935_4156.n5 a_3935_4156.t0 3.55417
R16964 a_3935_4156.t1 a_3935_4156.n5 3.32705
R16965 a_3935_4156.n4 a_3935_4156.t2 3.09022
R16966 a_3935_4156.n5 a_3935_4156.n4 1.2245
R16967 a_3935_4156.n1 a_3935_4156.n0 0.774747
R16968 a_3935_4156.n2 a_3935_4156.n1 0.774747
R16969 a_33216_1944.n10 a_33216_1944.t9 15.8415
R16970 a_33216_1944.n4 a_33216_1944.t13 15.8415
R16971 a_33216_1944.n5 a_33216_1944.t8 15.8415
R16972 a_33216_1944.n6 a_33216_1944.t12 15.8415
R16973 a_33216_1944.n7 a_33216_1944.t21 15.8415
R16974 a_33216_1944.n8 a_33216_1944.t23 15.8415
R16975 a_33216_1944.n9 a_33216_1944.t11 15.8415
R16976 a_33216_1944.n11 a_33216_1944.t22 15.8415
R16977 a_33216_1944.n10 a_33216_1944.t17 13.4447
R16978 a_33216_1944.n4 a_33216_1944.t20 13.4447
R16979 a_33216_1944.n5 a_33216_1944.t16 13.4447
R16980 a_33216_1944.n6 a_33216_1944.t19 13.4447
R16981 a_33216_1944.n7 a_33216_1944.t10 13.4447
R16982 a_33216_1944.n8 a_33216_1944.t15 13.4447
R16983 a_33216_1944.n9 a_33216_1944.t18 13.4447
R16984 a_33216_1944.n11 a_33216_1944.t14 13.4447
R16985 a_33216_1944.n5 a_33216_1944.n4 10.5449
R16986 a_33216_1944.n6 a_33216_1944.n5 10.5449
R16987 a_33216_1944.n7 a_33216_1944.n6 10.5449
R16988 a_33216_1944.n8 a_33216_1944.n7 10.5449
R16989 a_33216_1944.n9 a_33216_1944.n8 10.5449
R16990 a_33216_1944.n11 a_33216_1944.n9 10.5449
R16991 a_33216_1944.n11 a_33216_1944.n10 10.5449
R16992 a_33216_1944.n0 a_33216_1944.n3 7.22489
R16993 a_33216_1944.n0 a_33216_1944.n2 6.36702
R16994 a_33216_1944.n12 a_33216_1944.n0 3.56115
R16995 a_33216_1944.n0 a_33216_1944.n1 2.68463
R16996 a_33216_1944.n0 a_33216_1944.n11 2.37181
R16997 a_33216_1944.n1 a_33216_1944.t6 2.06607
R16998 a_33216_1944.t7 a_33216_1944.n12 2.06607
R16999 a_33216_1944.n2 a_33216_1944.t3 1.99806
R17000 a_33216_1944.n2 a_33216_1944.t1 1.99806
R17001 a_33216_1944.n3 a_33216_1944.t0 1.99806
R17002 a_33216_1944.n3 a_33216_1944.t2 1.99806
R17003 a_33216_1944.n1 a_33216_1944.t4 1.4923
R17004 a_33216_1944.n12 a_33216_1944.t5 1.4923
R17005 OUT[1] OUT[1].n14 21.4925
R17006 OUT[1].n3 OUT[1].n2 6.90733
R17007 OUT[1].n3 OUT[1].n1 6.3768
R17008 OUT[1].n12 OUT[1].n0 6.3768
R17009 OUT[1].n14 OUT[1].n13 6.3005
R17010 OUT[1].n9 OUT[1].n8 3.23472
R17011 OUT[1].n6 OUT[1].n5 3.21104
R17012 OUT[1].n9 OUT[1].n7 2.7042
R17013 OUT[1].n6 OUT[1].n4 2.7042
R17014 OUT[1].n7 OUT[1].t12 2.06607
R17015 OUT[1].n8 OUT[1].t11 2.06607
R17016 OUT[1].n5 OUT[1].t14 2.06607
R17017 OUT[1].n4 OUT[1].t8 2.06607
R17018 OUT[1].n13 OUT[1].t6 1.99806
R17019 OUT[1].n13 OUT[1].t3 1.99806
R17020 OUT[1].n2 OUT[1].t0 1.99806
R17021 OUT[1].n2 OUT[1].t4 1.99806
R17022 OUT[1].n1 OUT[1].t1 1.99806
R17023 OUT[1].n1 OUT[1].t7 1.99806
R17024 OUT[1].n0 OUT[1].t5 1.99806
R17025 OUT[1].n0 OUT[1].t2 1.99806
R17026 OUT[1].n7 OUT[1].t10 1.4923
R17027 OUT[1].n8 OUT[1].t15 1.4923
R17028 OUT[1].n5 OUT[1].t9 1.4923
R17029 OUT[1].n4 OUT[1].t13 1.4923
R17030 OUT[1].n14 OUT[1].n12 0.577837
R17031 OUT[1].n11 OUT[1].n3 0.189974
R17032 OUT[1].n10 OUT[1].n6 0.175763
R17033 OUT[1].n10 OUT[1].n9 0.166289
R17034 OUT[1].n12 OUT[1].n11 0.152079
R17035 OUT[1].n11 OUT[1].n10 0.145625
R17036 a_21772_n11428.n5 a_21772_n11428.t18 15.8415
R17037 a_21772_n11428.n6 a_21772_n11428.t21 15.8415
R17038 a_21772_n11428.n7 a_21772_n11428.t23 15.8415
R17039 a_21772_n11428.n8 a_21772_n11428.t19 15.8415
R17040 a_21772_n11428.n9 a_21772_n11428.t14 15.8415
R17041 a_21772_n11428.n10 a_21772_n11428.t17 15.8415
R17042 a_21772_n11428.n4 a_21772_n11428.t22 15.8415
R17043 a_21772_n11428.n11 a_21772_n11428.t20 15.8415
R17044 a_21772_n11428.n5 a_21772_n11428.t11 13.4447
R17045 a_21772_n11428.n6 a_21772_n11428.t8 13.4447
R17046 a_21772_n11428.n7 a_21772_n11428.t16 13.4447
R17047 a_21772_n11428.n8 a_21772_n11428.t12 13.4447
R17048 a_21772_n11428.n9 a_21772_n11428.t9 13.4447
R17049 a_21772_n11428.n10 a_21772_n11428.t10 13.4447
R17050 a_21772_n11428.n4 a_21772_n11428.t15 13.4447
R17051 a_21772_n11428.n11 a_21772_n11428.t13 13.4447
R17052 a_21772_n11428.n6 a_21772_n11428.n5 10.5449
R17053 a_21772_n11428.n7 a_21772_n11428.n6 10.5449
R17054 a_21772_n11428.n8 a_21772_n11428.n7 10.5449
R17055 a_21772_n11428.n9 a_21772_n11428.n8 10.5449
R17056 a_21772_n11428.n10 a_21772_n11428.n9 10.5449
R17057 a_21772_n11428.n11 a_21772_n11428.n4 10.5449
R17058 a_21772_n11428.n11 a_21772_n11428.n10 10.5449
R17059 a_21772_n11428.n0 a_21772_n11428.n3 7.22489
R17060 a_21772_n11428.n0 a_21772_n11428.n2 6.36702
R17061 a_21772_n11428.n12 a_21772_n11428.n0 3.56115
R17062 a_21772_n11428.n0 a_21772_n11428.n1 2.68463
R17063 a_21772_n11428.n0 a_21772_n11428.n11 2.37183
R17064 a_21772_n11428.n1 a_21772_n11428.t5 2.06607
R17065 a_21772_n11428.t7 a_21772_n11428.n12 2.06607
R17066 a_21772_n11428.n2 a_21772_n11428.t3 1.99806
R17067 a_21772_n11428.n2 a_21772_n11428.t2 1.99806
R17068 a_21772_n11428.n3 a_21772_n11428.t1 1.99806
R17069 a_21772_n11428.n3 a_21772_n11428.t0 1.99806
R17070 a_21772_n11428.n1 a_21772_n11428.t6 1.4923
R17071 a_21772_n11428.n12 a_21772_n11428.t4 1.4923
R17072 a_33496_n8222.n5 a_33496_n8222.t11 15.7685
R17073 a_33496_n8222.n6 a_33496_n8222.t21 15.7685
R17074 a_33496_n8222.n7 a_33496_n8222.t18 15.7685
R17075 a_33496_n8222.n8 a_33496_n8222.t9 15.7685
R17076 a_33496_n8222.n9 a_33496_n8222.t16 15.7685
R17077 a_33496_n8222.n10 a_33496_n8222.t15 15.7685
R17078 a_33496_n8222.n3 a_33496_n8222.t13 15.7685
R17079 a_33496_n8222.n4 a_33496_n8222.t20 15.7685
R17080 a_33496_n8222.n5 a_33496_n8222.t19 11.6197
R17081 a_33496_n8222.n6 a_33496_n8222.t22 11.6197
R17082 a_33496_n8222.n7 a_33496_n8222.t8 11.6197
R17083 a_33496_n8222.n8 a_33496_n8222.t10 11.6197
R17084 a_33496_n8222.n9 a_33496_n8222.t7 11.6197
R17085 a_33496_n8222.n10 a_33496_n8222.t17 11.6197
R17086 a_33496_n8222.n3 a_33496_n8222.t14 11.6197
R17087 a_33496_n8222.n4 a_33496_n8222.t12 11.6197
R17088 a_33496_n8222.n6 a_33496_n8222.n5 10.5449
R17089 a_33496_n8222.n7 a_33496_n8222.n6 10.5449
R17090 a_33496_n8222.n8 a_33496_n8222.n7 10.5449
R17091 a_33496_n8222.n9 a_33496_n8222.n8 10.5449
R17092 a_33496_n8222.n10 a_33496_n8222.n9 10.5449
R17093 a_33496_n8222.n4 a_33496_n8222.n3 10.5449
R17094 a_33496_n8222.n0 a_33496_n8222.t1 10.4819
R17095 a_33496_n8222.n11 a_33496_n8222.n10 8.41578
R17096 a_33496_n8222.n0 a_33496_n8222.n2 7.31398
R17097 a_33496_n8222.n12 a_33496_n8222.n0 6.25311
R17098 a_33496_n8222.n0 a_33496_n8222.n1 5.37659
R17099 a_33496_n8222.n2 a_33496_n8222.t0 4.04494
R17100 a_33496_n8222.n2 a_33496_n8222.t2 4.04494
R17101 a_33496_n8222.n1 a_33496_n8222.t3 3.07367
R17102 a_33496_n8222.n1 a_33496_n8222.t5 3.07367
R17103 a_33496_n8222.t6 a_33496_n8222.n12 3.07367
R17104 a_33496_n8222.n12 a_33496_n8222.t4 3.07367
R17105 a_33496_n8222.n0 a_33496_n8222.n11 2.93567
R17106 a_33496_n8222.n11 a_33496_n8222.n4 2.12967
R17107 a_31548_n10172.n17 a_31548_n10172.n16 25.5789
R17108 a_31548_n10172.n14 a_31548_n10172.n13 23.4189
R17109 a_31548_n10172.n12 a_31548_n10172.n11 23.2673
R17110 a_31548_n10172.n17 a_31548_n10172.n15 17.6873
R17111 a_31548_n10172.n12 a_31548_n10172.n10 17.6589
R17112 a_31548_n10172.n10 a_31548_n10172.t19 13.615
R17113 a_31548_n10172.n11 a_31548_n10172.t24 13.615
R17114 a_31548_n10172.n13 a_31548_n10172.t16 13.5542
R17115 a_31548_n10172.n15 a_31548_n10172.t18 13.5542
R17116 a_31548_n10172.n16 a_31548_n10172.t20 13.5542
R17117 a_31548_n10172.n13 a_31548_n10172.t25 12.4105
R17118 a_31548_n10172.n15 a_31548_n10172.t23 12.4105
R17119 a_31548_n10172.n16 a_31548_n10172.t21 12.4105
R17120 a_31548_n10172.n10 a_31548_n10172.t22 12.3375
R17121 a_31548_n10172.n11 a_31548_n10172.t17 12.3375
R17122 a_31548_n10172.n2 a_31548_n10172.n8 7.13263
R17123 a_31548_n10172.n0 a_31548_n10172.n6 7.13263
R17124 a_31548_n10172.n2 a_31548_n10172.n7 6.43746
R17125 a_31548_n10172.n0 a_31548_n10172.n5 6.43746
R17126 a_31548_n10172.n1 a_31548_n10172.n18 4.5005
R17127 a_31548_n10172.n18 a_31548_n10172.n17 4.3655
R17128 a_31548_n10172.n7 a_31548_n10172.t2 3.8098
R17129 a_31548_n10172.n7 a_31548_n10172.t7 3.8098
R17130 a_31548_n10172.n8 a_31548_n10172.t3 3.8098
R17131 a_31548_n10172.n8 a_31548_n10172.t4 3.8098
R17132 a_31548_n10172.n6 a_31548_n10172.t0 3.8098
R17133 a_31548_n10172.n6 a_31548_n10172.t1 3.8098
R17134 a_31548_n10172.n5 a_31548_n10172.t5 3.8098
R17135 a_31548_n10172.n5 a_31548_n10172.t6 3.8098
R17136 a_31548_n10172.n0 a_31548_n10172.n4 3.34593
R17137 a_31548_n10172.n1 a_31548_n10172.n9 2.94656
R17138 a_31548_n10172.n0 a_31548_n10172.n3 2.71593
R17139 a_31548_n10172.n19 a_31548_n10172.n0 2.71593
R17140 a_31548_n10172.n4 a_31548_n10172.t13 2.06607
R17141 a_31548_n10172.n4 a_31548_n10172.t9 2.06607
R17142 a_31548_n10172.n3 a_31548_n10172.t12 2.06607
R17143 a_31548_n10172.n3 a_31548_n10172.t11 2.06607
R17144 a_31548_n10172.n9 a_31548_n10172.t8 2.06607
R17145 a_31548_n10172.n9 a_31548_n10172.t14 2.06607
R17146 a_31548_n10172.t15 a_31548_n10172.n19 2.06607
R17147 a_31548_n10172.n19 a_31548_n10172.t10 2.06607
R17148 a_31548_n10172.n18 a_31548_n10172.n14 1.2155
R17149 a_31548_n10172.n14 a_31548_n10172.n12 1.0805
R17150 a_31548_n10172.n0 a_31548_n10172.n2 1.02848
R17151 a_31548_n10172.n0 a_31548_n10172.n1 0.745813
R17152 a_13501_n11816.n1 a_13501_n11816.t12 15.8618
R17153 a_13501_n11816.n0 a_13501_n11816.t13 15.8393
R17154 a_13501_n11816.n1 a_13501_n11816.t6 15.7537
R17155 a_13501_n11816.n0 a_13501_n11816.t5 15.7496
R17156 a_13501_n11816.n0 a_13501_n11816.n2 14.963
R17157 a_13501_n11816.n1 a_13501_n11816.n4 14.9583
R17158 a_13501_n11816.n1 a_13501_n11816.n8 14.9559
R17159 a_13501_n11816.n1 a_13501_n11816.n7 14.9547
R17160 a_13501_n11816.n0 a_13501_n11816.n3 14.7096
R17161 a_13501_n11816.n1 a_13501_n11816.n6 14.7035
R17162 a_13501_n11816.n1 a_13501_n11816.n5 14.7035
R17163 a_13501_n11816.n9 a_13501_n11816.n1 14.6941
R17164 a_13501_n11816.n6 a_13501_n11816.t8 0.6505
R17165 a_13501_n11816.n6 a_13501_n11816.t1 0.6505
R17166 a_13501_n11816.n5 a_13501_n11816.t0 0.6505
R17167 a_13501_n11816.n5 a_13501_n11816.t4 0.6505
R17168 a_13501_n11816.n3 a_13501_n11816.t3 0.6505
R17169 a_13501_n11816.n3 a_13501_n11816.t7 0.6505
R17170 a_13501_n11816.t9 a_13501_n11816.n9 0.6505
R17171 a_13501_n11816.n9 a_13501_n11816.t2 0.6505
R17172 a_13501_n11816.n8 a_13501_n11816.t19 0.5855
R17173 a_13501_n11816.n8 a_13501_n11816.t16 0.5855
R17174 a_13501_n11816.n7 a_13501_n11816.t10 0.5855
R17175 a_13501_n11816.n7 a_13501_n11816.t17 0.5855
R17176 a_13501_n11816.n4 a_13501_n11816.t18 0.5855
R17177 a_13501_n11816.n4 a_13501_n11816.t14 0.5855
R17178 a_13501_n11816.n2 a_13501_n11816.t15 0.5855
R17179 a_13501_n11816.n2 a_13501_n11816.t11 0.5855
R17180 a_13501_n11816.n1 a_13501_n11816.n0 0.158862
R17181 a_30732_332.n0 a_30732_332.t5 29.2005
R17182 a_30732_332.n2 a_30732_332.n0 27.5856
R17183 a_30732_332.t1 a_30732_332.n3 27.3145
R17184 a_30732_332.n1 a_30732_332.t2 19.7105
R17185 a_30732_332.n3 a_30732_332.t6 17.2528
R17186 a_30732_332.n1 a_30732_332.t7 13.3108
R17187 a_30732_332.t1 a_30732_332.t0 13.2903
R17188 a_30732_332.n2 a_30732_332.n1 13.1209
R17189 a_30732_332.n3 a_30732_332.t4 12.1672
R17190 a_30732_332.n0 a_30732_332.t3 12.1428
R17191 a_30732_332.t1 a_30732_332.n2 9.9005
R17192 a_21772_n452.n2 a_21772_n452.t8 15.8415
R17193 a_21772_n452.n3 a_21772_n452.t6 15.8415
R17194 a_21772_n452.n4 a_21772_n452.t9 15.8415
R17195 a_21772_n452.n5 a_21772_n452.t5 15.8415
R17196 a_21772_n452.n6 a_21772_n452.t15 15.8415
R17197 a_21772_n452.n7 a_21772_n452.t4 15.8415
R17198 a_21772_n452.n1 a_21772_n452.t7 15.8415
R17199 a_21772_n452.n0 a_21772_n452.t19 15.8415
R17200 a_21772_n452.n2 a_21772_n452.t12 13.4447
R17201 a_21772_n452.n3 a_21772_n452.t10 13.4447
R17202 a_21772_n452.n4 a_21772_n452.t17 13.4447
R17203 a_21772_n452.n5 a_21772_n452.t13 13.4447
R17204 a_21772_n452.n6 a_21772_n452.t11 13.4447
R17205 a_21772_n452.n7 a_21772_n452.t16 13.4447
R17206 a_21772_n452.n1 a_21772_n452.t18 13.4447
R17207 a_21772_n452.n0 a_21772_n452.t14 13.4447
R17208 a_21772_n452.n3 a_21772_n452.n2 10.5449
R17209 a_21772_n452.n4 a_21772_n452.n3 10.5449
R17210 a_21772_n452.n5 a_21772_n452.n4 10.5449
R17211 a_21772_n452.n6 a_21772_n452.n5 10.5449
R17212 a_21772_n452.n7 a_21772_n452.n6 10.5449
R17213 a_21772_n452.n0 a_21772_n452.n1 10.5449
R17214 a_21772_n452.n0 a_21772_n452.n7 10.5449
R17215 a_21772_n452.n0 a_21772_n452.t3 7.22489
R17216 a_21772_n452.n0 a_21772_n452.t1 7.12153
R17217 a_21772_n452.n0 a_21772_n452.t2 6.36702
R17218 a_21772_n452.t0 a_21772_n452.n0 5.62673
R17219 a_27259_804.n2 a_27259_804.n4 30.5295
R17220 a_27259_804.n0 a_27259_804.n3 29.6258
R17221 a_27259_804.n9 a_27259_804.n8 19.4672
R17222 a_27259_804.n10 a_27259_804.n7 19.4672
R17223 a_27259_804.n6 a_27259_804.t14 19.0535
R17224 a_27259_804.n3 a_27259_804.t13 18.9805
R17225 a_27259_804.n1 a_27259_804.t19 18.7737
R17226 a_27259_804.n4 a_27259_804.t4 18.6885
R17227 a_27259_804.n1 a_27259_804.n6 16.5048
R17228 a_27259_804.n8 a_27259_804.t11 16.4255
R17229 a_27259_804.n8 a_27259_804.t9 16.3282
R17230 a_27259_804.n9 a_27259_804.t7 15.9875
R17231 a_27259_804.n7 a_27259_804.t15 15.9875
R17232 a_27259_804.n10 a_27259_804.t17 15.9875
R17233 a_27259_804.n5 a_27259_804.t12 15.3305
R17234 a_27259_804.n5 a_27259_804.t6 15.0872
R17235 a_27259_804.n6 a_27259_804.t3 14.7952
R17236 a_27259_804.n9 a_27259_804.t18 14.7222
R17237 a_27259_804.n7 a_27259_804.t8 14.7222
R17238 a_27259_804.n10 a_27259_804.t10 14.7222
R17239 a_27259_804.n2 a_27259_804.n1 14.6546
R17240 a_27259_804.n0 a_27259_804.n2 13.5005
R17241 a_27259_804.n1 a_27259_804.t16 13.4447
R17242 a_27259_804.n2 a_27259_804.n5 12.5111
R17243 a_27259_804.n4 a_27259_804.t5 11.8752
R17244 a_27259_804.n3 a_27259_804.t2 11.4372
R17245 a_27259_804.n10 a_27259_804.n9 10.5449
R17246 a_27259_804.t1 a_27259_804.n0 9.42921
R17247 a_27259_804.n2 a_27259_804.n10 7.43285
R17248 a_27259_804.n0 a_27259_804.t0 7.34176
R17249 a_25612_n878.n4 a_25612_n878.n2 21.5722
R17250 a_25612_n878.n5 a_25612_n878.n4 19.3505
R17251 a_25612_n878.n1 a_25612_n878.t4 18.9805
R17252 a_25612_n878.n3 a_25612_n878.t2 18.6885
R17253 a_25612_n878.n2 a_25612_n878.t6 17.484
R17254 a_25612_n878.n5 a_25612_n878.n1 16.6646
R17255 a_25612_n878.n4 a_25612_n878.n3 13.4107
R17256 a_25612_n878.n3 a_25612_n878.t7 11.9603
R17257 a_25612_n878.n2 a_25612_n878.t5 11.863
R17258 a_25612_n878.n1 a_25612_n878.t3 11.4372
R17259 a_25612_n878.n0 a_25612_n878.t1 8.31075
R17260 a_25612_n878.n0 a_25612_n878.n5 6.0755
R17261 a_25612_n878.t0 a_25612_n878.n0 5.13976
R17262 a_28519_n10160.n2 a_28519_n10160.t5 19.4185
R17263 a_28519_n10160.n1 a_28519_n10160.t2 19.2725
R17264 a_28519_n10160.n0 a_28519_n10160.t8 17.5205
R17265 a_28519_n10160.n5 a_28519_n10160.n4 17.2446
R17266 a_28519_n10160.n4 a_28519_n10160.t9 17.119
R17267 a_28519_n10160.n3 a_28519_n10160.n0 15.0932
R17268 a_28519_n10160.n3 a_28519_n10160.n2 13.5355
R17269 a_28519_n10160.n5 a_28519_n10160.n3 12.9605
R17270 a_28519_n10160.n4 a_28519_n10160.t6 12.7147
R17271 a_28519_n10160.n3 a_28519_n10160.n1 12.7017
R17272 a_28519_n10160.t1 a_28519_n10160.n5 11.7005
R17273 a_28519_n10160.n2 a_28519_n10160.t3 11.6683
R17274 a_28519_n10160.n0 a_28519_n10160.t4 11.5588
R17275 a_28519_n10160.n1 a_28519_n10160.t7 10.9505
R17276 a_28519_n10160.t1 a_28519_n10160.t0 8.30886
R17277 a_22220_690.n8 a_22220_690.n6 34.7486
R17278 a_22220_690.n10 a_22220_690.n2 31.1405
R17279 a_22220_690.n2 a_22220_690.n1 23.2478
R17280 a_22220_690.n1 a_22220_690.n3 20.0181
R17281 a_22220_690.n4 a_22220_690.t16 18.9805
R17282 a_22220_690.n9 a_22220_690.t2 18.6885
R17283 a_22220_690.n2 a_22220_690.n5 17.6508
R17284 a_22220_690.n6 a_22220_690.t8 17.484
R17285 a_22220_690.n5 a_22220_690.t7 15.4522
R17286 a_22220_690.n5 a_22220_690.t9 15.1115
R17287 a_22220_690.n1 a_22220_690.n4 13.9658
R17288 a_22220_690.n10 a_22220_690.n9 12.7042
R17289 a_22220_690.n9 a_22220_690.t17 11.8752
R17290 a_22220_690.n6 a_22220_690.t12 11.863
R17291 a_22220_690.t1 a_22220_690.n12 11.5205
R17292 a_22220_690.n4 a_22220_690.t14 11.4372
R17293 a_22220_690.n12 a_22220_690.n10 10.6205
R17294 a_22220_690.n2 a_22220_690.n8 10.0355
R17295 a_22220_690.n12 a_22220_690.n11 9.0005
R17296 a_22220_690.n1 a_22220_690.n0 9.0005
R17297 a_22220_690.t1 a_22220_690.t0 8.60215
R17298 a_22220_690.n0 a_22220_690.t10 6.71423
R17299 a_22220_690.n11 a_22220_690.t4 6.56378
R17300 a_22220_690.n7 a_22220_690.t6 6.3005
R17301 a_22220_690.n3 a_22220_690.t13 6.3005
R17302 a_22220_690.n7 a_22220_690.t15 5.6196
R17303 a_22220_690.n3 a_22220_690.t11 5.6196
R17304 a_22220_690.n11 a_22220_690.t3 5.35632
R17305 a_22220_690.n0 a_22220_690.t5 5.20587
R17306 a_22220_690.n8 a_22220_690.n7 4.53811
R17307 OUT[3] OUT[3].n14 20.8003
R17308 OUT[3].n9 OUT[3].n8 6.90733
R17309 OUT[3].n6 OUT[3].n5 6.89497
R17310 OUT[3].n9 OUT[3].n7 6.3768
R17311 OUT[3].n6 OUT[3].n4 6.3768
R17312 OUT[3].n3 OUT[3].n2 3.23472
R17313 OUT[3].n3 OUT[3].n1 2.7042
R17314 OUT[3].n12 OUT[3].n0 2.7042
R17315 OUT[3].n14 OUT[3].n13 2.6005
R17316 OUT[3].n13 OUT[3].t15 2.06607
R17317 OUT[3].n2 OUT[3].t12 2.06607
R17318 OUT[3].n1 OUT[3].t8 2.06607
R17319 OUT[3].n0 OUT[3].t13 2.06607
R17320 OUT[3].n7 OUT[3].t1 1.99806
R17321 OUT[3].n7 OUT[3].t7 1.99806
R17322 OUT[3].n8 OUT[3].t5 1.99806
R17323 OUT[3].n8 OUT[3].t3 1.99806
R17324 OUT[3].n5 OUT[3].t2 1.99806
R17325 OUT[3].n5 OUT[3].t0 1.99806
R17326 OUT[3].n4 OUT[3].t6 1.99806
R17327 OUT[3].n4 OUT[3].t4 1.99806
R17328 OUT[3].n13 OUT[3].t9 1.4923
R17329 OUT[3].n2 OUT[3].t10 1.4923
R17330 OUT[3].n1 OUT[3].t14 1.4923
R17331 OUT[3].n0 OUT[3].t11 1.4923
R17332 OUT[3].n14 OUT[3].n12 0.601315
R17333 OUT[3].n10 OUT[3].n9 0.189974
R17334 OUT[3].n12 OUT[3].n11 0.175763
R17335 OUT[3].n11 OUT[3].n3 0.166289
R17336 OUT[3].n10 OUT[3].n6 0.152079
R17337 OUT[3].n11 OUT[3].n10 0.145625
R17338 a_21692_n5111.n3 a_21692_n5111.n2 31.0955
R17339 a_21692_n5111.n2 a_21692_n5111.n0 30.1287
R17340 a_21692_n5111.n0 a_21692_n5111.t3 19.7105
R17341 a_21692_n5111.n1 a_21692_n5111.t4 19.7105
R17342 a_21692_n5111.n0 a_21692_n5111.t2 13.3108
R17343 a_21692_n5111.n1 a_21692_n5111.t5 13.3108
R17344 a_21692_n5111.n3 a_21692_n5111.t0 9.61569
R17345 a_21692_n5111.n2 a_21692_n5111.n1 8.7537
R17346 a_21692_n5111.t1 a_21692_n5111.n3 4.52215
R17347 a_13501_n22528.n1 a_13501_n22528.t3 15.8618
R17348 a_13501_n22528.n0 a_13501_n22528.t2 15.8393
R17349 a_13501_n22528.n1 a_13501_n22528.t12 15.7537
R17350 a_13501_n22528.n0 a_13501_n22528.t11 15.7496
R17351 a_13501_n22528.n0 a_13501_n22528.n2 14.963
R17352 a_13501_n22528.n1 a_13501_n22528.n4 14.9583
R17353 a_13501_n22528.n1 a_13501_n22528.n8 14.9559
R17354 a_13501_n22528.n1 a_13501_n22528.n7 14.9547
R17355 a_13501_n22528.n0 a_13501_n22528.n3 14.7096
R17356 a_13501_n22528.n1 a_13501_n22528.n6 14.7035
R17357 a_13501_n22528.n1 a_13501_n22528.n5 14.7035
R17358 a_13501_n22528.n9 a_13501_n22528.n1 14.6941
R17359 a_13501_n22528.n6 a_13501_n22528.t14 0.6505
R17360 a_13501_n22528.n6 a_13501_n22528.t17 0.6505
R17361 a_13501_n22528.n5 a_13501_n22528.t16 0.6505
R17362 a_13501_n22528.n5 a_13501_n22528.t10 0.6505
R17363 a_13501_n22528.n3 a_13501_n22528.t19 0.6505
R17364 a_13501_n22528.n3 a_13501_n22528.t13 0.6505
R17365 a_13501_n22528.n9 a_13501_n22528.t15 0.6505
R17366 a_13501_n22528.t18 a_13501_n22528.n9 0.6505
R17367 a_13501_n22528.n8 a_13501_n22528.t6 0.5855
R17368 a_13501_n22528.n8 a_13501_n22528.t9 0.5855
R17369 a_13501_n22528.n7 a_13501_n22528.t5 0.5855
R17370 a_13501_n22528.n7 a_13501_n22528.t8 0.5855
R17371 a_13501_n22528.n4 a_13501_n22528.t7 0.5855
R17372 a_13501_n22528.n4 a_13501_n22528.t1 0.5855
R17373 a_13501_n22528.n2 a_13501_n22528.t0 0.5855
R17374 a_13501_n22528.n2 a_13501_n22528.t4 0.5855
R17375 a_13501_n22528.n1 a_13501_n22528.n0 0.158862
R17376 a_24481_761.t80 a_24481_761.t89 274.176
R17377 a_24481_761.t33 a_24481_761.t29 254.709
R17378 a_24481_761.t46 a_24481_761.t31 254.709
R17379 a_24481_761.t93 a_24481_761.t87 254.709
R17380 a_24481_761.t8 a_24481_761.t22 254.709
R17381 a_24481_761.t68 a_24481_761.t35 254.709
R17382 a_24481_761.t70 a_24481_761.t28 254.709
R17383 a_24481_761.t12 a_24481_761.t61 254.709
R17384 a_24481_761.t71 a_24481_761.t51 254.709
R17385 a_24481_761.t15 a_24481_761.t94 254.709
R17386 a_24481_761.t73 a_24481_761.t77 254.709
R17387 a_24481_761.t39 a_24481_761.t30 254.709
R17388 a_24481_761.t82 a_24481_761.t45 211.846
R17389 a_24481_761.n44 a_24481_761.t74 31.6987
R17390 a_24481_761.n36 a_24481_761.t72 31.4493
R17391 a_24481_761.n24 a_24481_761.t86 31.4493
R17392 a_24481_761.n16 a_24481_761.t84 31.4493
R17393 a_24481_761.n20 a_24481_761.t58 31.4493
R17394 a_24481_761.n17 a_24481_761.t56 31.4493
R17395 a_24481_761.n33 a_24481_761.t11 31.4493
R17396 a_24481_761.n27 a_24481_761.t54 31.4493
R17397 a_24481_761.n28 a_24481_761.t49 31.4493
R17398 a_24481_761.n39 a_24481_761.t38 31.4493
R17399 a_24481_761.n42 a_24481_761.t41 31.4493
R17400 a_24481_761.n34 a_24481_761.t18 29.8433
R17401 a_24481_761.n38 a_24481_761.t13 29.8433
R17402 a_24481_761.n30 a_24481_761.n28 25.7363
R17403 a_24481_761.t29 a_24481_761.t62 23.7012
R17404 a_24481_761.t31 a_24481_761.t66 23.7012
R17405 a_24481_761.t87 a_24481_761.t14 23.7012
R17406 a_24481_761.t89 a_24481_761.t27 23.7012
R17407 a_24481_761.t22 a_24481_761.t67 23.7012
R17408 a_24481_761.t35 a_24481_761.t90 23.7012
R17409 a_24481_761.t28 a_24481_761.t60 23.7012
R17410 a_24481_761.t61 a_24481_761.t21 23.7012
R17411 a_24481_761.t51 a_24481_761.t81 23.7012
R17412 a_24481_761.t94 a_24481_761.t9 23.7012
R17413 a_24481_761.t77 a_24481_761.t64 23.7012
R17414 a_24481_761.t30 a_24481_761.t32 23.7012
R17415 a_24481_761.t45 a_24481_761.t50 23.4396
R17416 a_24481_761.n5 a_24481_761.n34 21.7345
R17417 a_24481_761.n46 a_24481_761.n43 20.5205
R17418 a_24481_761.n0 a_24481_761.n2 19.3259
R17419 a_24481_761.n43 a_24481_761.n42 18.815
R17420 a_24481_761.n45 a_24481_761.t26 18.6885
R17421 a_24481_761.n2 a_24481_761.t88 18.6885
R17422 a_24481_761.n44 a_24481_761.t23 18.6885
R17423 a_24481_761.n3 a_24481_761.n24 17.0963
R17424 a_24481_761.n40 a_24481_761.n38 16.9138
R17425 a_24481_761.n19 a_24481_761.n17 15.08
R17426 a_24481_761.n10 a_24481_761.n40 14.5805
R17427 a_24481_761.n18 a_24481_761.t78 14.2998
R17428 a_24481_761.n18 a_24481_761.t82 13.8705
R17429 a_24481_761.n1 a_24481_761.n20 13.86
R17430 a_24481_761.n40 a_24481_761.n39 13.7663
R17431 a_24481_761.n7 a_24481_761.n27 13.46
R17432 a_24481_761.n11 a_24481_761.n16 12.92
R17433 a_24481_761.n7 a_24481_761.n33 12.5963
R17434 a_24481_761.n19 a_24481_761.n18 12.5159
R17435 a_24481_761.n37 a_24481_761.n36 12.5038
R17436 a_24481_761.n11 a_24481_761.n22 11.8355
R17437 a_24481_761.n22 a_24481_761.n19 11.2955
R17438 a_24481_761.n45 a_24481_761.t40 11.1938
R17439 a_24481_761.n2 a_24481_761.t20 11.1938
R17440 a_24481_761.n44 a_24481_761.t37 11.1938
R17441 a_24481_761.n32 a_24481_761.n31 10.9731
R17442 a_24481_761.n2 a_24481_761.n45 10.5449
R17443 a_24481_761.n2 a_24481_761.n44 10.5449
R17444 a_24481_761.n3 a_24481_761.n15 10.2981
R17445 a_24481_761.n10 a_24481_761.n4 10.0805
R17446 a_24481_761.n4 a_24481_761.n13 9.75811
R17447 a_24481_761.n0 a_24481_761.t25 9.70587
R17448 a_24481_761.n4 a_24481_761.n14 9.5405
R17449 a_24481_761.n8 a_24481_761.n46 9.5405
R17450 a_24481_761.n22 a_24481_761.n1 9.2705
R17451 a_24481_761.n6 a_24481_761.n3 8.3705
R17452 a_24481_761.n4 a_24481_761.n37 7.9205
R17453 a_24481_761.n7 a_24481_761.n32 7.7405
R17454 a_24481_761.n32 a_24481_761.n30 7.5605
R17455 a_24481_761.n3 a_24481_761.n11 7.2905
R17456 a_24481_761.n5 a_24481_761.n7 7.2005
R17457 a_24481_761.n8 a_24481_761.t7 7.13263
R17458 a_24481_761.n8 a_24481_761.t6 7.13263
R17459 a_24481_761.n6 a_24481_761.n5 6.9755
R17460 a_24481_761.n7 a_24481_761.n26 6.92311
R17461 a_24481_761.n36 a_24481_761.t33 6.79462
R17462 a_24481_761.n24 a_24481_761.t46 6.79462
R17463 a_24481_761.n16 a_24481_761.t93 6.79462
R17464 a_24481_761.n17 a_24481_761.t8 6.79462
R17465 a_24481_761.n34 a_24481_761.t68 6.79462
R17466 a_24481_761.n33 a_24481_761.t70 6.79462
R17467 a_24481_761.n27 a_24481_761.t12 6.79462
R17468 a_24481_761.n28 a_24481_761.t71 6.79462
R17469 a_24481_761.n38 a_24481_761.t15 6.79462
R17470 a_24481_761.n39 a_24481_761.t73 6.79462
R17471 a_24481_761.n42 a_24481_761.t39 6.79462
R17472 a_24481_761.n0 a_24481_761.t91 6.71423
R17473 a_24481_761.n12 a_24481_761.t47 6.71423
R17474 a_24481_761.n21 a_24481_761.t92 6.71423
R17475 a_24481_761.n1 a_24481_761.t17 6.71423
R17476 a_24481_761.n9 a_24481_761.t75 6.56378
R17477 a_24481_761.n8 a_24481_761.t4 6.43746
R17478 a_24481_761.n8 a_24481_761.t5 6.43746
R17479 a_24481_761.n14 a_24481_761.t19 6.41334
R17480 a_24481_761.n35 a_24481_761.t76 6.3005
R17481 a_24481_761.n25 a_24481_761.t43 6.3005
R17482 a_24481_761.n15 a_24481_761.t63 6.3005
R17483 a_24481_761.n23 a_24481_761.t83 6.3005
R17484 a_24481_761.n26 a_24481_761.t52 6.3005
R17485 a_24481_761.n29 a_24481_761.t79 6.3005
R17486 a_24481_761.n31 a_24481_761.t55 6.3005
R17487 a_24481_761.n13 a_24481_761.t85 6.3005
R17488 a_24481_761.n20 a_24481_761.t80 6.0198
R17489 a_24481_761.n35 a_24481_761.t34 5.6196
R17490 a_24481_761.n25 a_24481_761.t24 5.6196
R17491 a_24481_761.n15 a_24481_761.t44 5.6196
R17492 a_24481_761.n23 a_24481_761.t57 5.6196
R17493 a_24481_761.n26 a_24481_761.t16 5.6196
R17494 a_24481_761.n29 a_24481_761.t53 5.6196
R17495 a_24481_761.n31 a_24481_761.t65 5.6196
R17496 a_24481_761.n13 a_24481_761.t59 5.6196
R17497 a_24481_761.n43 a_24481_761.n41 5.5805
R17498 a_24481_761.n10 a_24481_761.n9 5.5805
R17499 a_24481_761.n41 a_24481_761.n12 5.5355
R17500 a_24481_761.n14 a_24481_761.t10 5.50677
R17501 a_24481_761.n46 a_24481_761.n0 5.4005
R17502 a_24481_761.n9 a_24481_761.t69 5.35632
R17503 a_24481_761.t0 a_24481_761.n8 5.27673
R17504 a_24481_761.n1 a_24481_761.n21 5.2205
R17505 a_24481_761.n11 a_24481_761.n23 5.21311
R17506 a_24481_761.n12 a_24481_761.t42 5.20587
R17507 a_24481_761.n21 a_24481_761.t36 5.20587
R17508 a_24481_761.n1 a_24481_761.t48 5.20587
R17509 a_24481_761.n41 a_24481_761.n10 5.1755
R17510 a_24481_761.n8 a_24481_761.t1 4.85463
R17511 a_24481_761.n8 a_24481_761.t3 4.78151
R17512 a_24481_761.n8 a_24481_761.t2 4.78151
R17513 a_24481_761.n37 a_24481_761.n6 4.6355
R17514 a_24481_761.n6 a_24481_761.n35 4.53811
R17515 a_24481_761.n6 a_24481_761.n25 4.53811
R17516 a_24481_761.n30 a_24481_761.n29 4.53811
R17517 a_26328_n6654.n5 a_26328_n6654.t20 15.7685
R17518 a_26328_n6654.n6 a_26328_n6654.t13 15.7685
R17519 a_26328_n6654.n7 a_26328_n6654.t21 15.7685
R17520 a_26328_n6654.n8 a_26328_n6654.t16 15.7685
R17521 a_26328_n6654.n9 a_26328_n6654.t9 15.7685
R17522 a_26328_n6654.n10 a_26328_n6654.t19 15.7685
R17523 a_26328_n6654.n3 a_26328_n6654.t10 15.7685
R17524 a_26328_n6654.n4 a_26328_n6654.t11 15.7685
R17525 a_26328_n6654.n5 a_26328_n6654.t7 11.6197
R17526 a_26328_n6654.n6 a_26328_n6654.t22 11.6197
R17527 a_26328_n6654.n7 a_26328_n6654.t8 11.6197
R17528 a_26328_n6654.n8 a_26328_n6654.t12 11.6197
R17529 a_26328_n6654.n9 a_26328_n6654.t14 11.6197
R17530 a_26328_n6654.n10 a_26328_n6654.t17 11.6197
R17531 a_26328_n6654.n3 a_26328_n6654.t18 11.6197
R17532 a_26328_n6654.n4 a_26328_n6654.t15 11.6197
R17533 a_26328_n6654.n6 a_26328_n6654.n5 10.5449
R17534 a_26328_n6654.n7 a_26328_n6654.n6 10.5449
R17535 a_26328_n6654.n8 a_26328_n6654.n7 10.5449
R17536 a_26328_n6654.n9 a_26328_n6654.n8 10.5449
R17537 a_26328_n6654.n10 a_26328_n6654.n9 10.5449
R17538 a_26328_n6654.n4 a_26328_n6654.n3 10.5449
R17539 a_26328_n6654.n0 a_26328_n6654.t1 10.4819
R17540 a_26328_n6654.n11 a_26328_n6654.n10 8.41578
R17541 a_26328_n6654.n0 a_26328_n6654.n2 7.31398
R17542 a_26328_n6654.n0 a_26328_n6654.n1 6.25311
R17543 a_26328_n6654.n12 a_26328_n6654.n0 5.37659
R17544 a_26328_n6654.n2 a_26328_n6654.t2 4.04494
R17545 a_26328_n6654.n2 a_26328_n6654.t0 4.04494
R17546 a_26328_n6654.n1 a_26328_n6654.t4 3.07367
R17547 a_26328_n6654.n1 a_26328_n6654.t3 3.07367
R17548 a_26328_n6654.t6 a_26328_n6654.n12 3.07367
R17549 a_26328_n6654.n12 a_26328_n6654.t5 3.07367
R17550 a_26328_n6654.n0 a_26328_n6654.n11 2.93567
R17551 a_26328_n6654.n11 a_26328_n6654.n4 2.12967
R17552 a_21692_n13308.n1 a_21692_n13308.n22 22.0955
R17553 a_21692_n13308.n13 a_21692_n13308.n12 18.3789
R17554 a_21692_n13308.n11 a_21692_n13308.n10 17.1473
R17555 a_21692_n13308.n9 a_21692_n13308.n7 15.9489
R17556 a_21692_n13308.n10 a_21692_n13308.t22 13.615
R17557 a_21692_n13308.n8 a_21692_n13308.t18 13.615
R17558 a_21692_n13308.n7 a_21692_n13308.t21 13.615
R17559 a_21692_n13308.n6 a_21692_n13308.t17 13.5542
R17560 a_21692_n13308.n20 a_21692_n13308.t19 13.5542
R17561 a_21692_n13308.n18 a_21692_n13308.t28 13.5542
R17562 a_21692_n13308.n16 a_21692_n13308.t29 13.5542
R17563 a_21692_n13308.n12 a_21692_n13308.t30 13.5542
R17564 a_21692_n13308.n14 a_21692_n13308.t27 13.5542
R17565 a_21692_n13308.n15 a_21692_n13308.n14 12.7989
R17566 a_21692_n13308.n11 a_21692_n13308.n9 12.7805
R17567 a_21692_n13308.n17 a_21692_n13308.n16 12.6473
R17568 a_21692_n13308.n22 a_21692_n13308.n6 12.6189
R17569 a_21692_n13308.n21 a_21692_n13308.n20 12.6189
R17570 a_21692_n13308.n19 a_21692_n13308.n18 12.6189
R17571 a_21692_n13308.n9 a_21692_n13308.n8 12.5147
R17572 a_21692_n13308.n6 a_21692_n13308.t26 12.4105
R17573 a_21692_n13308.n20 a_21692_n13308.t33 12.4105
R17574 a_21692_n13308.n18 a_21692_n13308.t32 12.4105
R17575 a_21692_n13308.n16 a_21692_n13308.t16 12.4105
R17576 a_21692_n13308.n12 a_21692_n13308.t24 12.4105
R17577 a_21692_n13308.n14 a_21692_n13308.t31 12.4105
R17578 a_21692_n13308.n10 a_21692_n13308.t25 12.3375
R17579 a_21692_n13308.n8 a_21692_n13308.t23 12.3375
R17580 a_21692_n13308.n7 a_21692_n13308.t20 12.3375
R17581 a_21692_n13308.n15 a_21692_n13308.n13 7.6955
R17582 a_21692_n13308.n0 a_21692_n13308.n26 7.13263
R17583 a_21692_n13308.n0 a_21692_n13308.n24 7.13263
R17584 a_21692_n13308.n0 a_21692_n13308.n25 6.43746
R17585 a_21692_n13308.n0 a_21692_n13308.n23 6.43746
R17586 a_21692_n13308.n13 a_21692_n13308.n11 5.4005
R17587 a_21692_n13308.n25 a_21692_n13308.t2 3.8098
R17588 a_21692_n13308.n25 a_21692_n13308.t4 3.8098
R17589 a_21692_n13308.n26 a_21692_n13308.t1 3.8098
R17590 a_21692_n13308.n26 a_21692_n13308.t3 3.8098
R17591 a_21692_n13308.n24 a_21692_n13308.t0 3.8098
R17592 a_21692_n13308.n24 a_21692_n13308.t7 3.8098
R17593 a_21692_n13308.n23 a_21692_n13308.t5 3.8098
R17594 a_21692_n13308.n23 a_21692_n13308.t6 3.8098
R17595 a_21692_n13308.n2 a_21692_n13308.n3 3.34593
R17596 a_21692_n13308.n22 a_21692_n13308.n21 3.1055
R17597 a_21692_n13308.n1 a_21692_n13308.n5 3.10406
R17598 a_21692_n13308.n2 a_21692_n13308.n4 2.71593
R17599 a_21692_n13308.n27 a_21692_n13308.n2 2.71593
R17600 a_21692_n13308.n19 a_21692_n13308.n17 2.6555
R17601 a_21692_n13308.n21 a_21692_n13308.n19 2.5205
R17602 a_21692_n13308.n17 a_21692_n13308.n15 2.4305
R17603 a_21692_n13308.n4 a_21692_n13308.t11 2.06607
R17604 a_21692_n13308.n4 a_21692_n13308.t8 2.06607
R17605 a_21692_n13308.n5 a_21692_n13308.t12 2.06607
R17606 a_21692_n13308.n5 a_21692_n13308.t9 2.06607
R17607 a_21692_n13308.n3 a_21692_n13308.t14 2.06607
R17608 a_21692_n13308.n3 a_21692_n13308.t13 2.06607
R17609 a_21692_n13308.n27 a_21692_n13308.t10 2.06607
R17610 a_21692_n13308.t15 a_21692_n13308.n27 2.06607
R17611 a_21692_n13308.n2 a_21692_n13308.n0 0.851294
R17612 a_21692_n13308.n2 a_21692_n13308.n1 0.7655
R17613 a_30452_n5156.n11 a_30452_n5156.n10 30.4701
R17614 a_30452_n5156.n7 a_30452_n5156.n6 30.4701
R17615 a_30452_n5156.n14 a_30452_n5156.n13 23.0405
R17616 a_30452_n5156.n13 a_30452_n5156.n0 19.6624
R17617 a_30452_n5156.n11 a_30452_n5156.t8 18.9805
R17618 a_30452_n5156.n10 a_30452_n5156.t3 18.9805
R17619 a_30452_n5156.n6 a_30452_n5156.t14 18.9805
R17620 a_30452_n5156.n7 a_30452_n5156.t6 18.9805
R17621 a_30452_n5156.n3 a_30452_n5156.t10 15.8415
R17622 a_30452_n5156.n2 a_30452_n5156.t9 15.8415
R17623 a_30452_n5156.n3 a_30452_n5156.t4 13.4447
R17624 a_30452_n5156.n2 a_30452_n5156.t5 13.4447
R17625 a_30452_n5156.n12 a_30452_n5156.t13 10.5612
R17626 a_30452_n5156.n9 a_30452_n5156.t12 10.5612
R17627 a_30452_n5156.n5 a_30452_n5156.t7 10.5612
R17628 a_30452_n5156.n8 a_30452_n5156.t11 10.5612
R17629 a_30452_n5156.n0 a_30452_n5156.n12 9.70845
R17630 a_30452_n5156.n0 a_30452_n5156.n5 8.54637
R17631 a_30452_n5156.n0 a_30452_n5156.n8 8.0005
R17632 a_30452_n5156.n9 a_30452_n5156.n0 8.0005
R17633 a_30452_n5156.n13 a_30452_n5156.n4 7.30054
R17634 a_30452_n5156.n14 a_30452_n5156.n1 7.08733
R17635 a_30452_n5156.n4 a_30452_n5156.n2 6.388
R17636 a_30452_n5156.n4 a_30452_n5156.n3 4.76578
R17637 a_30452_n5156.n12 a_30452_n5156.n11 4.2345
R17638 a_30452_n5156.n10 a_30452_n5156.n9 4.2345
R17639 a_30452_n5156.n6 a_30452_n5156.n5 4.2345
R17640 a_30452_n5156.n8 a_30452_n5156.n7 4.2345
R17641 a_30452_n5156.n1 a_30452_n5156.t0 3.37782
R17642 a_30452_n5156.n1 a_30452_n5156.t1 3.37782
R17643 a_30452_n5156.t2 a_30452_n5156.n14 2.78525
R17644 a_28736_n4633.n15 a_28736_n4633.n14 28.3769
R17645 a_28736_n4633.n2 a_28736_n4633.t22 20.9945
R17646 a_28736_n4633.n14 a_28736_n4633.t23 17.7395
R17647 a_28736_n4633.n2 a_28736_n4633.t21 17.2189
R17648 a_28736_n4633.n13 a_28736_n4633.t25 16.1822
R17649 a_28736_n4633.n13 a_28736_n4633.t20 14.0165
R17650 a_28736_n4633.n14 a_28736_n4633.t24 12.6782
R17651 a_28736_n4633.n2 a_28736_n4633.n13 8.39556
R17652 a_28736_n4633.n5 a_28736_n4633.n3 8.0692
R17653 a_28736_n4633.n15 a_28736_n4633.n2 7.33492
R17654 a_28736_n4633.n5 a_28736_n4633.n4 6.3005
R17655 a_28736_n4633.n0 a_28736_n4633.n12 6.03444
R17656 a_28736_n4633.n0 a_28736_n4633.n15 5.7605
R17657 a_28736_n4633.n1 a_28736_n4633.n6 5.3668
R17658 a_28736_n4633.n1 a_28736_n4633.n7 5.3668
R17659 a_28736_n4633.n1 a_28736_n4633.n8 5.3668
R17660 a_28736_n4633.n0 a_28736_n4633.n9 5.3668
R17661 a_28736_n4633.n0 a_28736_n4633.n10 5.3668
R17662 a_28736_n4633.n0 a_28736_n4633.n11 5.3668
R17663 a_28736_n4633.n17 a_28736_n4633.n16 5.3668
R17664 a_28736_n4633.n3 a_28736_n4633.t16 3.6883
R17665 a_28736_n4633.n3 a_28736_n4633.t15 3.6883
R17666 a_28736_n4633.n4 a_28736_n4633.t14 3.6883
R17667 a_28736_n4633.n4 a_28736_n4633.t17 3.6883
R17668 a_28736_n4633.n16 a_28736_n4633.n1 2.29141
R17669 a_28736_n4633.n6 a_28736_n4633.t12 2.15435
R17670 a_28736_n4633.n6 a_28736_n4633.t0 2.15435
R17671 a_28736_n4633.n7 a_28736_n4633.t1 2.15435
R17672 a_28736_n4633.n7 a_28736_n4633.t13 2.15435
R17673 a_28736_n4633.n8 a_28736_n4633.t11 2.15435
R17674 a_28736_n4633.n8 a_28736_n4633.t2 2.15435
R17675 a_28736_n4633.n9 a_28736_n4633.t8 2.15435
R17676 a_28736_n4633.n9 a_28736_n4633.t5 2.15435
R17677 a_28736_n4633.n10 a_28736_n4633.t4 2.15435
R17678 a_28736_n4633.n10 a_28736_n4633.t9 2.15435
R17679 a_28736_n4633.n11 a_28736_n4633.t7 2.15435
R17680 a_28736_n4633.n11 a_28736_n4633.t6 2.15435
R17681 a_28736_n4633.n12 a_28736_n4633.t19 2.15435
R17682 a_28736_n4633.n12 a_28736_n4633.t18 2.15435
R17683 a_28736_n4633.t3 a_28736_n4633.n17 2.15435
R17684 a_28736_n4633.n17 a_28736_n4633.t10 2.15435
R17685 a_28736_n4633.n1 a_28736_n4633.n0 2.00341
R17686 a_28736_n4633.n16 a_28736_n4633.n5 1.64833
R17687 a_35456_n4628.n8 a_35456_n4628.t22 15.7685
R17688 a_35456_n4628.n9 a_35456_n4628.t19 15.7685
R17689 a_35456_n4628.n2 a_35456_n4628.t13 15.7685
R17690 a_35456_n4628.n3 a_35456_n4628.t18 15.7685
R17691 a_35456_n4628.n4 a_35456_n4628.t11 15.7685
R17692 a_35456_n4628.n5 a_35456_n4628.t12 15.7685
R17693 a_35456_n4628.n6 a_35456_n4628.t20 15.7685
R17694 a_35456_n4628.n7 a_35456_n4628.t14 15.7685
R17695 a_35456_n4628.n8 a_35456_n4628.t21 11.6197
R17696 a_35456_n4628.n9 a_35456_n4628.t7 11.6197
R17697 a_35456_n4628.n2 a_35456_n4628.t17 11.6197
R17698 a_35456_n4628.n3 a_35456_n4628.t15 11.6197
R17699 a_35456_n4628.n4 a_35456_n4628.t16 11.6197
R17700 a_35456_n4628.n5 a_35456_n4628.t9 11.6197
R17701 a_35456_n4628.n6 a_35456_n4628.t8 11.6197
R17702 a_35456_n4628.n7 a_35456_n4628.t10 11.6197
R17703 a_35456_n4628.n9 a_35456_n4628.n8 10.5449
R17704 a_35456_n4628.n3 a_35456_n4628.n2 10.5449
R17705 a_35456_n4628.n4 a_35456_n4628.n3 10.5449
R17706 a_35456_n4628.n5 a_35456_n4628.n4 10.5449
R17707 a_35456_n4628.n6 a_35456_n4628.n5 10.5449
R17708 a_35456_n4628.n7 a_35456_n4628.n6 10.5449
R17709 a_35456_n4628.n0 a_35456_n4628.t0 10.4819
R17710 a_35456_n4628.n10 a_35456_n4628.n7 8.41578
R17711 a_35456_n4628.n0 a_35456_n4628.n1 7.31398
R17712 a_35456_n4628.n0 a_35456_n4628.n11 6.25311
R17713 a_35456_n4628.n12 a_35456_n4628.n0 5.37659
R17714 a_35456_n4628.n1 a_35456_n4628.t2 4.04494
R17715 a_35456_n4628.n1 a_35456_n4628.t1 4.04494
R17716 a_35456_n4628.n11 a_35456_n4628.t5 3.07367
R17717 a_35456_n4628.n11 a_35456_n4628.t3 3.07367
R17718 a_35456_n4628.n12 a_35456_n4628.t4 3.07367
R17719 a_35456_n4628.t6 a_35456_n4628.n12 3.07367
R17720 a_35456_n4628.n0 a_35456_n4628.n10 2.93567
R17721 a_35456_n4628.n10 a_35456_n4628.n9 2.12967
R17722 a_32108_n2332.n14 a_32108_n2332.n13 26.6589
R17723 a_32108_n2332.n10 a_32108_n2332.n9 17.1473
R17724 a_32108_n2332.n0 a_32108_n2332.n16 15.9755
R17725 a_32108_n2332.n8 a_32108_n2332.n6 14.0139
R17726 a_32108_n2332.n11 a_32108_n2332.t24 13.615
R17727 a_32108_n2332.n9 a_32108_n2332.t20 13.615
R17728 a_32108_n2332.n7 a_32108_n2332.t18 13.615
R17729 a_32108_n2332.n15 a_32108_n2332.t25 13.5542
R17730 a_32108_n2332.n6 a_32108_n2332.t21 13.5542
R17731 a_32108_n2332.n13 a_32108_n2332.t26 13.5542
R17732 a_32108_n2332.n16 a_32108_n2332.n15 12.6473
R17733 a_32108_n2332.n8 a_32108_n2332.n7 12.6473
R17734 a_32108_n2332.n12 a_32108_n2332.n11 12.6189
R17735 a_32108_n2332.n15 a_32108_n2332.t19 12.4105
R17736 a_32108_n2332.n6 a_32108_n2332.t23 12.4105
R17737 a_32108_n2332.n13 a_32108_n2332.t27 12.4105
R17738 a_32108_n2332.n11 a_32108_n2332.t22 12.3375
R17739 a_32108_n2332.n9 a_32108_n2332.t16 12.3375
R17740 a_32108_n2332.n7 a_32108_n2332.t17 12.3375
R17741 a_32108_n2332.n10 a_32108_n2332.n8 11.1605
R17742 a_32108_n2332.n12 a_32108_n2332.n10 9.7205
R17743 a_32108_n2332.n1 a_32108_n2332.n20 7.13263
R17744 a_32108_n2332.n2 a_32108_n2332.n18 7.13263
R17745 a_32108_n2332.n1 a_32108_n2332.n19 6.43746
R17746 a_32108_n2332.n2 a_32108_n2332.n17 6.43746
R17747 a_32108_n2332.n19 a_32108_n2332.t2 3.8098
R17748 a_32108_n2332.n19 a_32108_n2332.t5 3.8098
R17749 a_32108_n2332.n20 a_32108_n2332.t1 3.8098
R17750 a_32108_n2332.n20 a_32108_n2332.t3 3.8098
R17751 a_32108_n2332.n18 a_32108_n2332.t7 3.8098
R17752 a_32108_n2332.n18 a_32108_n2332.t0 3.8098
R17753 a_32108_n2332.n17 a_32108_n2332.t6 3.8098
R17754 a_32108_n2332.n17 a_32108_n2332.t4 3.8098
R17755 a_32108_n2332.n14 a_32108_n2332.n12 3.7805
R17756 a_32108_n2332.n0 a_32108_n2332.n3 3.34593
R17757 a_32108_n2332.n0 a_32108_n2332.n5 2.80031
R17758 a_32108_n2332.n16 a_32108_n2332.n14 2.7455
R17759 a_32108_n2332.n0 a_32108_n2332.n4 2.71593
R17760 a_32108_n2332.n21 a_32108_n2332.n0 2.71593
R17761 a_32108_n2332.n4 a_32108_n2332.t9 2.06607
R17762 a_32108_n2332.n4 a_32108_n2332.t12 2.06607
R17763 a_32108_n2332.n5 a_32108_n2332.t10 2.06607
R17764 a_32108_n2332.n5 a_32108_n2332.t8 2.06607
R17765 a_32108_n2332.n3 a_32108_n2332.t13 2.06607
R17766 a_32108_n2332.n3 a_32108_n2332.t11 2.06607
R17767 a_32108_n2332.t15 a_32108_n2332.n21 2.06607
R17768 a_32108_n2332.n21 a_32108_n2332.t14 2.06607
R17769 a_32108_n2332.n0 a_32108_n2332.n1 1.3428
R17770 a_32108_n2332.n1 a_32108_n2332.n2 0.577741
R17771 a_25940_n17606.n20 a_25940_n17606.n0 21.9155
R17772 a_25940_n17606.n2 a_25940_n17606.n17 19.1705
R17773 a_25940_n17606.n18 a_25940_n17606.t5 17.8003
R17774 a_25940_n17606.n16 a_25940_n17606.t8 17.7395
R17775 a_25940_n17606.n11 a_25940_n17606.t3 17.7395
R17776 a_25940_n17606.n7 a_25940_n17606.t2 17.7395
R17777 a_25940_n17606.n6 a_25940_n17606.t6 17.7395
R17778 a_25940_n17606.n0 a_25940_n17606.n2 16.5155
R17779 a_25940_n17606.n1 a_25940_n17606.n4 16.2005
R17780 a_25940_n17606.n3 a_25940_n17606.t9 16.1822
R17781 a_25940_n17606.n3 a_25940_n17606.t7 14.8925
R17782 a_25940_n17606.n18 a_25940_n17606.t13 14.8195
R17783 a_25940_n17606.n17 a_25940_n17606.n16 13.7969
R17784 a_25940_n17606.n2 a_25940_n17606.n18 13.4692
R17785 a_25940_n17606.n0 a_25940_n17606.n3 12.7152
R17786 a_25940_n17606.n16 a_25940_n17606.t19 12.6782
R17787 a_25940_n17606.n11 a_25940_n17606.t15 12.6782
R17788 a_25940_n17606.n7 a_25940_n17606.t22 12.6782
R17789 a_25940_n17606.n6 a_25940_n17606.t11 12.6782
R17790 a_25940_n17606.n10 a_25940_n17606.n8 11.5205
R17791 a_25940_n17606.n8 a_25940_n17606.n7 8.92214
R17792 a_25940_n17606.n13 a_25940_n17606.n11 8.84694
R17793 a_25940_n17606.n1 a_25940_n17606.n6 8.57694
R17794 a_25940_n17606.n0 a_25940_n17606.n19 6.83311
R17795 a_25940_n17606.n5 a_25940_n17606.t25 6.71423
R17796 a_25940_n17606.n20 a_25940_n17606.t0 6.69707
R17797 a_25940_n17606.n17 a_25940_n17606.n15 6.4805
R17798 a_25940_n17606.n4 a_25940_n17606.t14 6.41334
R17799 a_25940_n17606.n14 a_25940_n17606.t21 6.3005
R17800 a_25940_n17606.n12 a_25940_n17606.t12 6.3005
R17801 a_25940_n17606.n9 a_25940_n17606.t17 6.3005
R17802 a_25940_n17606.n19 a_25940_n17606.t16 6.3005
R17803 a_25940_n17606.n14 a_25940_n17606.t20 5.6196
R17804 a_25940_n17606.n12 a_25940_n17606.t10 5.6196
R17805 a_25940_n17606.n9 a_25940_n17606.t18 5.6196
R17806 a_25940_n17606.n19 a_25940_n17606.t24 5.6196
R17807 a_25940_n17606.n4 a_25940_n17606.t23 5.50677
R17808 a_25940_n17606.n5 a_25940_n17606.t4 5.20587
R17809 a_25940_n17606.n13 a_25940_n17606.n12 5.07811
R17810 a_25940_n17606.n8 a_25940_n17606.n1 4.8155
R17811 a_25940_n17606.n10 a_25940_n17606.n9 4.71811
R17812 a_25940_n17606.n15 a_25940_n17606.n14 4.53811
R17813 a_25940_n17606.n1 a_25940_n17606.n5 4.5005
R17814 a_25940_n17606.n2 a_25940_n17606.n10 4.0505
R17815 a_25940_n17606.t1 a_25940_n17606.n20 3.0803
R17816 a_25940_n17606.n15 a_25940_n17606.n13 2.4755
R17817 a_22140_n6694.n14 a_22140_n6694.n0 22.7711
R17818 a_22140_n6694.n8 a_22140_n6694.t2 18.9805
R17819 a_22140_n6694.n3 a_22140_n6694.t8 18.6885
R17820 a_22140_n6694.n5 a_22140_n6694.t3 18.6885
R17821 a_22140_n6694.n14 a_22140_n6694.n13 16.0205
R17822 a_22140_n6694.n0 a_22140_n6694.t17 15.3305
R17823 a_22140_n6694.n0 a_22140_n6694.t13 15.148
R17824 a_22140_n6694.n4 a_22140_n6694.n3 13.2661
R17825 a_22140_n6694.n10 a_22140_n6694.n8 12.7538
R17826 a_22140_n6694.n3 a_22140_n6694.t4 11.9603
R17827 a_22140_n6694.n5 a_22140_n6694.t15 11.9603
R17828 a_22140_n6694.n8 a_22140_n6694.t5 11.4372
R17829 a_22140_n6694.n7 a_22140_n6694.n1 11.3405
R17830 a_22140_n6694.n11 a_22140_n6694.n7 11.2505
R17831 a_22140_n6694.n13 a_22140_n6694.n12 10.8005
R17832 a_22140_n6694.n4 a_22140_n6694.n2 10.6205
R17833 a_22140_n6694.n11 a_22140_n6694.n10 10.5755
R17834 a_22140_n6694.t1 a_22140_n6694.n14 10.4405
R17835 a_22140_n6694.n6 a_22140_n6694.n5 8.85295
R17836 a_22140_n6694.n6 a_22140_n6694.n4 8.5955
R17837 a_22140_n6694.t1 a_22140_n6694.t0 8.30886
R17838 a_22140_n6694.n10 a_22140_n6694.n9 7.55311
R17839 a_22140_n6694.n7 a_22140_n6694.n6 6.9755
R17840 a_22140_n6694.n12 a_22140_n6694.t10 6.71423
R17841 a_22140_n6694.n1 a_22140_n6694.t16 6.71423
R17842 a_22140_n6694.n2 a_22140_n6694.t6 6.56378
R17843 a_22140_n6694.n9 a_22140_n6694.t14 6.3005
R17844 a_22140_n6694.n9 a_22140_n6694.t9 5.6196
R17845 a_22140_n6694.n13 a_22140_n6694.n11 5.5805
R17846 a_22140_n6694.n2 a_22140_n6694.t7 5.35632
R17847 a_22140_n6694.n12 a_22140_n6694.t11 5.20587
R17848 a_22140_n6694.n1 a_22140_n6694.t12 5.20587
R17849 a_22672_n2214.n1 a_22672_n2214.n0 43.2816
R17850 a_22672_n2214.n0 a_22672_n2214.t3 29.2005
R17851 a_22672_n2214.n0 a_22672_n2214.t4 12.1428
R17852 a_22672_n2214.n1 a_22672_n2214.t2 6.58175
R17853 a_22672_n2214.t2 a_22672_n2214.t0 5.92991
R17854 a_22672_n2214.t1 a_22672_n2214.n1 5.69912
R17855 a_29444_n4328.n3 a_29444_n4328.n2 46.4036
R17856 a_29444_n4328.n2 a_29444_n4328.t9 17.484
R17857 a_29444_n4328.n1 a_29444_n4328.t6 17.3015
R17858 a_29444_n4328.n3 a_29444_n4328.n1 17.1981
R17859 a_29444_n4328.n2 a_29444_n4328.t7 11.863
R17860 a_29444_n4328.n1 a_29444_n4328.t8 10.6463
R17861 a_29444_n4328.n0 a_29444_n4328.t0 8.32963
R17862 a_29444_n4328.n0 a_29444_n4328.t4 7.90366
R17863 a_29444_n4328.n0 a_29444_n4328.t5 7.44983
R17864 a_29444_n4328.n0 a_29444_n4328.n3 6.33857
R17865 a_29444_n4328.t1 a_29444_n4328.n0 5.2005
R17866 a_29444_n4328.n0 a_29444_n4328.t2 5.2005
R17867 a_29444_n4328.n0 a_29444_n4328.t3 5.2005
R17868 a_29900_760.n7 a_29900_760.n3 22.6805
R17869 a_29900_760.n0 a_29900_760.t5 20.9945
R17870 a_29900_760.n2 a_29900_760.t7 20.9945
R17871 a_29900_760.n1 a_29900_760.t13 20.9945
R17872 a_29900_760.n3 a_29900_760.t3 20.9945
R17873 a_29900_760.n4 a_29900_760.n2 19.9355
R17874 a_29900_760.n4 a_29900_760.n7 17.6405
R17875 a_29900_760.n0 a_29900_760.t11 17.2633
R17876 a_29900_760.n1 a_29900_760.t8 17.2633
R17877 a_29900_760.n3 a_29900_760.t14 17.0442
R17878 a_29900_760.n2 a_29900_760.t15 16.9182
R17879 a_29900_760.n9 a_29900_760.t9 16.1822
R17880 a_29900_760.n8 a_29900_760.t6 16.1822
R17881 a_29900_760.n6 a_29900_760.t16 16.1822
R17882 a_29900_760.n5 a_29900_760.t12 16.1822
R17883 a_29900_760.n9 a_29900_760.t4 14.0165
R17884 a_29900_760.n8 a_29900_760.t2 14.0165
R17885 a_29900_760.n6 a_29900_760.t10 14.0165
R17886 a_29900_760.n5 a_29900_760.t17 14.0165
R17887 a_29900_760.n2 a_29900_760.n8 8.74067
R17888 a_29900_760.n3 a_29900_760.n5 8.61467
R17889 a_29900_760.n0 a_29900_760.n9 8.04725
R17890 a_29900_760.n1 a_29900_760.n6 8.04725
R17891 a_29900_760.n10 a_29900_760.t0 7.02633
R17892 a_29900_760.n10 a_29900_760.n4 5.8955
R17893 a_29900_760.n4 a_29900_760.n0 5.02881
R17894 a_29900_760.n7 a_29900_760.n1 4.84881
R17895 a_29900_760.t1 a_29900_760.n10 2.74964
R17896 a_11023_n4162.n19 a_11023_n4162.t37 56.0276
R17897 a_11023_n4162.n10 a_11023_n4162.t36 56.019
R17898 a_11023_n4162.n12 a_11023_n4162.t26 55.9719
R17899 a_11023_n4162.n6 a_11023_n4162.t35 55.9719
R17900 a_11023_n4162.n14 a_11023_n4162.t31 55.9719
R17901 a_11023_n4162.n5 a_11023_n4162.t23 55.9719
R17902 a_11023_n4162.n16 a_11023_n4162.t33 55.9719
R17903 a_11023_n4162.n4 a_11023_n4162.t28 55.9719
R17904 a_11023_n4162.n17 a_11023_n4162.t39 55.9719
R17905 a_11023_n4162.n2 a_11023_n4162.t34 55.9719
R17906 a_11023_n4162.n20 a_11023_n4162.t30 55.9719
R17907 a_11023_n4162.n10 a_11023_n4162.t25 55.9719
R17908 a_11023_n4162.n10 a_11023_n4162.t21 55.9719
R17909 a_11023_n4162.n9 a_11023_n4162.t38 55.9719
R17910 a_11023_n4162.n9 a_11023_n4162.t27 55.9719
R17911 a_11023_n4162.n7 a_11023_n4162.t22 55.9719
R17912 a_11023_n4162.n7 a_11023_n4162.t32 55.9719
R17913 a_11023_n4162.n8 a_11023_n4162.t24 55.9719
R17914 a_11023_n4162.n8 a_11023_n4162.t20 55.9719
R17915 a_11023_n4162.n25 a_11023_n4162.t29 55.9719
R17916 a_11023_n4162.n12 a_11023_n4162.n11 0.0590857
R17917 a_11023_n4162.n22 a_11023_n4162.n21 4.5005
R17918 a_11023_n4162.n23 a_11023_n4162.n2 4.5005
R17919 a_11023_n4162.n17 a_11023_n4162.n24 4.5005
R17920 a_11023_n4162.n3 a_11023_n4162.n0 4.5005
R17921 a_11023_n4162.n1 a_11023_n4162.n4 4.5005
R17922 a_11023_n4162.n16 a_11023_n4162.n15 4.5005
R17923 a_11023_n4162.n31 a_11023_n4162.n30 4.5005
R17924 a_11023_n4162.n29 a_11023_n4162.n5 4.5005
R17925 a_11023_n4162.n14 a_11023_n4162.n13 4.5005
R17926 a_11023_n4162.n28 a_11023_n4162.n27 4.5005
R17927 a_11023_n4162.n26 a_11023_n4162.n6 4.5005
R17928 a_11023_n4162.n37 a_11023_n4162.n36 3.87048
R17929 a_11023_n4162.n37 a_11023_n4162.n35 3.68704
R17930 a_11023_n4162.n38 a_11023_n4162.n34 3.68704
R17931 a_11023_n4162.n39 a_11023_n4162.n33 3.68704
R17932 a_11023_n4162.n40 a_11023_n4162.n32 3.68704
R17933 a_11023_n4162.n48 a_11023_n4162.n18 3.53719
R17934 a_11023_n4162.n43 a_11023_n4162.n42 3.37808
R17935 a_11023_n4162.n45 a_11023_n4162.n44 3.37808
R17936 a_11023_n4162.n47 a_11023_n4162.n46 3.37808
R17937 a_11023_n4162.n49 a_11023_n4162.n48 3.37783
R17938 a_11023_n4162.n41 a_11023_n4162.n1 1.89107
R17939 a_11023_n4162.n22 a_11023_n4162.n19 1.15666
R17940 a_11023_n4162.n42 a_11023_n4162.t16 0.6505
R17941 a_11023_n4162.n42 a_11023_n4162.t14 0.6505
R17942 a_11023_n4162.n44 a_11023_n4162.t13 0.6505
R17943 a_11023_n4162.n44 a_11023_n4162.t10 0.6505
R17944 a_11023_n4162.n46 a_11023_n4162.t12 0.6505
R17945 a_11023_n4162.n46 a_11023_n4162.t18 0.6505
R17946 a_11023_n4162.n18 a_11023_n4162.t17 0.6505
R17947 a_11023_n4162.n18 a_11023_n4162.t11 0.6505
R17948 a_11023_n4162.t19 a_11023_n4162.n49 0.6505
R17949 a_11023_n4162.n49 a_11023_n4162.t15 0.6505
R17950 a_11023_n4162.n36 a_11023_n4162.t7 0.5855
R17951 a_11023_n4162.n36 a_11023_n4162.t1 0.5855
R17952 a_11023_n4162.n35 a_11023_n4162.t9 0.5855
R17953 a_11023_n4162.n35 a_11023_n4162.t5 0.5855
R17954 a_11023_n4162.n34 a_11023_n4162.t2 0.5855
R17955 a_11023_n4162.n34 a_11023_n4162.t8 0.5855
R17956 a_11023_n4162.n33 a_11023_n4162.t3 0.5855
R17957 a_11023_n4162.n33 a_11023_n4162.t0 0.5855
R17958 a_11023_n4162.n32 a_11023_n4162.t6 0.5855
R17959 a_11023_n4162.n32 a_11023_n4162.t4 0.5855
R17960 a_11023_n4162.n41 a_11023_n4162.n40 0.41138
R17961 a_11023_n4162.n43 a_11023_n4162.n41 0.373278
R17962 a_11023_n4162.n38 a_11023_n4162.n37 0.183939
R17963 a_11023_n4162.n39 a_11023_n4162.n38 0.183939
R17964 a_11023_n4162.n40 a_11023_n4162.n39 0.183939
R17965 a_11023_n4162.n48 a_11023_n4162.n47 0.159616
R17966 a_11023_n4162.n47 a_11023_n4162.n45 0.159616
R17967 a_11023_n4162.n45 a_11023_n4162.n43 0.159616
R17968 a_11023_n4162.n20 a_11023_n4162.n19 0.121859
R17969 a_11023_n4162.n21 a_11023_n4162.n20 0.11975
R17970 a_11023_n4162.n17 a_11023_n4162.n2 0.11975
R17971 a_11023_n4162.n4 a_11023_n4162.n16 0.11975
R17972 a_11023_n4162.n5 a_11023_n4162.n14 0.11975
R17973 a_11023_n4162.n6 a_11023_n4162.n12 0.11975
R17974 a_11023_n4162.n23 a_11023_n4162.n22 0.11975
R17975 a_11023_n4162.n24 a_11023_n4162.n23 0.11975
R17976 a_11023_n4162.n24 a_11023_n4162.n0 0.11975
R17977 a_11023_n4162.n1 a_11023_n4162.n15 0.11975
R17978 a_11023_n4162.n30 a_11023_n4162.n15 0.11975
R17979 a_11023_n4162.n30 a_11023_n4162.n29 0.11975
R17980 a_11023_n4162.n29 a_11023_n4162.n13 0.11975
R17981 a_11023_n4162.n27 a_11023_n4162.n13 0.11975
R17982 a_11023_n4162.n27 a_11023_n4162.n26 0.11975
R17983 a_11023_n4162.n26 a_11023_n4162.n11 2.37025
R17984 a_11023_n4162.n3 a_11023_n4162.n17 0.11975
R17985 a_11023_n4162.n16 a_11023_n4162.n31 0.11975
R17986 a_11023_n4162.n14 a_11023_n4162.n28 0.11975
R17987 a_11023_n4162.n11 a_11023_n4162.n25 1.35571
R17988 a_11023_n4162.n28 a_11023_n4162.n6 0.11975
R17989 a_11023_n4162.n31 a_11023_n4162.n5 0.11975
R17990 a_11023_n4162.n4 a_11023_n4162.n3 0.11975
R17991 a_11023_n4162.n21 a_11023_n4162.n2 0.11975
R17992 a_11023_n4162.n1 a_11023_n4162.n0 0.11975
R17993 a_11023_n4162.n9 a_11023_n4162.n10 0.0946176
R17994 a_11023_n4162.n7 a_11023_n4162.n9 0.0946176
R17995 a_11023_n4162.n8 a_11023_n4162.n7 0.0946176
R17996 a_11023_n4162.n25 a_11023_n4162.n8 0.0946176
R17997 a_11087_n20850.n40 a_11087_n20850.n39 318.031
R17998 a_11087_n20850.n33 a_11087_n20850.n32 76.5005
R17999 a_11087_n20850.n11 a_11087_n20850.n36 60.7605
R18000 a_11087_n20850.n32 a_11087_n20850.n17 58.5005
R18001 a_11087_n20850.n35 a_11087_n20850.n17 38.4755
R18002 a_11087_n20850.n36 a_11087_n20850.n35 38.0255
R18003 a_11087_n20850.n22 a_11087_n20850.t29 10.553
R18004 a_11087_n20850.n40 a_11087_n20850.t0 10.4369
R18005 a_11087_n20850.n41 a_11087_n20850.t14 10.4369
R18006 a_11087_n20850.n42 a_11087_n20850.t9 10.4308
R18007 a_11087_n20850.n43 a_11087_n20850.t11 10.4308
R18008 a_11087_n20850.n44 a_11087_n20850.t5 10.4308
R18009 a_11087_n20850.n22 a_11087_n20850.t21 10.4156
R18010 a_11087_n20850.n24 a_11087_n20850.t25 10.4129
R18011 a_11087_n20850.n25 a_11087_n20850.t26 10.4121
R18012 a_11087_n20850.n23 a_11087_n20850.t28 10.4121
R18013 a_11087_n20850.n49 a_11087_n20850.t10 10.357
R18014 a_11087_n20850.n46 a_11087_n20850.t16 10.2004
R18015 a_11087_n20850.n48 a_11087_n20850.t13 10.2004
R18016 a_11087_n20850.n47 a_11087_n20850.t18 10.198
R18017 a_11087_n20850.t7 a_11087_n20850.n49 10.1921
R18018 a_11087_n20850.n38 a_11087_n20850.n37 5.94277
R18019 a_11087_n20850.t33 a_11087_n20850.n21 1.49319
R18020 a_11087_n20850.n33 a_11087_n20850.n21 60.7744
R18021 a_11087_n20850.n37 a_11087_n20850.n6 4.52686
R18022 a_11087_n20850.n11 a_11087_n20850.n10 4.5005
R18023 a_11087_n20850.n5 a_11087_n20850.n27 4.52686
R18024 a_11087_n20850.n13 a_11087_n20850.n12 4.5005
R18025 a_11087_n20850.n34 a_11087_n20850.n16 4.52686
R18026 a_11087_n20850.n18 a_11087_n20850.n14 4.5005
R18027 a_11087_n20850.n7 a_11087_n20850.n31 4.52686
R18028 a_11087_n20850.n30 a_11087_n20850.n19 4.5005
R18029 a_11087_n20850.n29 a_11087_n20850.n9 4.52686
R18030 a_11087_n20850.n28 a_11087_n20850.n20 4.5005
R18031 a_11087_n20850.t37 a_11087_n20850.n2 1.13765
R18032 a_11087_n20850.t32 a_11087_n20850.n1 0.251795
R18033 a_11087_n20850.n0 a_11087_n20850.n38 3.14437
R18034 a_11087_n20850.n26 a_11087_n20850.n4 3.85832
R18035 a_11087_n20850.n11 a_11087_n20850.n6 0.0273431
R18036 a_11087_n20850.n5 a_11087_n20850.n13 0.0273431
R18037 a_11087_n20850.n18 a_11087_n20850.n16 0.0273431
R18038 a_11087_n20850.n19 a_11087_n20850.n7 0.0273431
R18039 a_11087_n20850.n20 a_11087_n20850.n9 0.0273431
R18040 a_11087_n20850.n36 a_11087_n20850.n13 2.26055
R18041 a_11087_n20850.n18 a_11087_n20850.n17 2.26055
R18042 a_11087_n20850.n32 a_11087_n20850.n19 2.26055
R18043 a_11087_n20850.n33 a_11087_n20850.n20 2.26055
R18044 a_11087_n20850.n30 a_11087_n20850.n29 1.83512
R18045 a_11087_n20850.n2 a_11087_n20850.n1 3.4891
R18046 a_11087_n20850.n39 a_11087_n20850.n0 2.30525
R18047 a_11087_n20850.n27 a_11087_n20850.n10 1.37358
R18048 a_11087_n20850.n31 a_11087_n20850.n14 1.37358
R18049 a_11087_n20850.n28 a_11087_n20850.n21 3.65519
R18050 a_11087_n20850.n1 a_11087_n20850.n39 31.6166
R18051 a_11087_n20850.n26 a_11087_n20850.n2 6.23969
R18052 a_11087_n20850.t38 a_11087_n20850.t31 1.56538
R18053 a_11087_n20850.n26 a_11087_n20850.t40 1.2147
R18054 a_11087_n20850.n38 a_11087_n20850.t39 1.0799
R18055 a_11087_n20850.t36 a_11087_n20850.t41 0.9605
R18056 a_11087_n20850.t36 a_11087_n20850.n3 0.0276952
R18057 a_11087_n20850.n35 a_11087_n20850.n34 0.923577
R18058 a_11087_n20850.n35 a_11087_n20850.n12 0.912038
R18059 a_11087_n20850.n46 a_11087_n20850.n45 0.773592
R18060 a_11087_n20850.t16 a_11087_n20850.t8 0.6505
R18061 a_11087_n20850.t18 a_11087_n20850.t3 0.6505
R18062 a_11087_n20850.t13 a_11087_n20850.t4 0.6505
R18063 a_11087_n20850.t10 a_11087_n20850.t15 0.6505
R18064 a_11087_n20850.t1 a_11087_n20850.t7 0.6505
R18065 a_11087_n20850.t26 a_11087_n20850.t20 0.5855
R18066 a_11087_n20850.t25 a_11087_n20850.t23 0.5855
R18067 a_11087_n20850.t28 a_11087_n20850.t22 0.5855
R18068 a_11087_n20850.t21 a_11087_n20850.t24 0.5855
R18069 a_11087_n20850.t29 a_11087_n20850.t27 0.5855
R18070 a_11087_n20850.t0 a_11087_n20850.t12 0.5855
R18071 a_11087_n20850.t14 a_11087_n20850.t6 0.5855
R18072 a_11087_n20850.t9 a_11087_n20850.t2 0.5855
R18073 a_11087_n20850.t11 a_11087_n20850.t17 0.5855
R18074 a_11087_n20850.t5 a_11087_n20850.t19 0.5855
R18075 a_11087_n20850.t31 a_11087_n20850.n0 1.10549
R18076 a_11087_n20850.n15 a_11087_n20850.t34 0.484786
R18077 a_11087_n20850.n45 a_11087_n20850.n25 0.365893
R18078 a_11087_n20850.t34 a_11087_n20850.n6 1.47948
R18079 a_11087_n20850.t34 a_11087_n20850.n5 1.45162
R18080 a_11087_n20850.n16 a_11087_n20850.n15 1.45162
R18081 a_11087_n20850.n8 a_11087_n20850.n7 1.45162
R18082 a_11087_n20850.t33 a_11087_n20850.n9 1.45162
R18083 a_11087_n20850.n45 a_11087_n20850.n44 0.297718
R18084 a_11087_n20850.n41 a_11087_n20850.n40 0.1615
R18085 a_11087_n20850.n47 a_11087_n20850.n46 0.161
R18086 a_11087_n20850.n44 a_11087_n20850.n43 0.1605
R18087 a_11087_n20850.n43 a_11087_n20850.n42 0.1605
R18088 a_11087_n20850.n49 a_11087_n20850.n48 0.1605
R18089 a_11087_n20850.n48 a_11087_n20850.n47 0.1605
R18090 a_11087_n20850.n42 a_11087_n20850.n41 0.1585
R18091 a_11087_n20850.n25 a_11087_n20850.n24 0.139126
R18092 a_11087_n20850.n23 a_11087_n20850.n22 0.136566
R18093 a_11087_n20850.n24 a_11087_n20850.n23 0.13486
R18094 a_11087_n20850.n37 a_11087_n20850.n10 0.127423
R18095 a_11087_n20850.n27 a_11087_n20850.n12 0.127423
R18096 a_11087_n20850.n34 a_11087_n20850.n14 0.127423
R18097 a_11087_n20850.n31 a_11087_n20850.n30 0.127423
R18098 a_11087_n20850.n29 a_11087_n20850.n28 0.127423
R18099 a_11087_n20850.n8 a_11087_n20850.t35 0.0708125
R18100 a_11087_n20850.n4 a_11087_n20850.t41 0.0343063
R18101 a_11087_n20850.n3 a_11087_n20850.t30 1.08464
R18102 a_11087_n20850.n8 a_11087_n20850.t33 0.512643
R18103 a_11087_n20850.n15 a_11087_n20850.n8 0.0562143
R18104 a_11087_n20850.n4 a_11087_n20850.n3 1.0109
R18105 a_11087_n20850.t32 a_11087_n20850.t37 0.996929
R18106 a_30192_n15304.n9 a_30192_n15304.t13 15.7685
R18107 a_30192_n15304.n10 a_30192_n15304.t7 15.7685
R18108 a_30192_n15304.n3 a_30192_n15304.t8 15.7685
R18109 a_30192_n15304.n4 a_30192_n15304.t10 15.7685
R18110 a_30192_n15304.n5 a_30192_n15304.t11 15.7685
R18111 a_30192_n15304.n6 a_30192_n15304.t9 15.7685
R18112 a_30192_n15304.n7 a_30192_n15304.t20 15.7685
R18113 a_30192_n15304.n8 a_30192_n15304.t12 15.7685
R18114 a_30192_n15304.n9 a_30192_n15304.t22 11.6197
R18115 a_30192_n15304.n10 a_30192_n15304.t17 11.6197
R18116 a_30192_n15304.n3 a_30192_n15304.t18 11.6197
R18117 a_30192_n15304.n4 a_30192_n15304.t16 11.6197
R18118 a_30192_n15304.n5 a_30192_n15304.t21 11.6197
R18119 a_30192_n15304.n6 a_30192_n15304.t15 11.6197
R18120 a_30192_n15304.n7 a_30192_n15304.t14 11.6197
R18121 a_30192_n15304.n8 a_30192_n15304.t19 11.6197
R18122 a_30192_n15304.n10 a_30192_n15304.n9 10.5449
R18123 a_30192_n15304.n4 a_30192_n15304.n3 10.5449
R18124 a_30192_n15304.n5 a_30192_n15304.n4 10.5449
R18125 a_30192_n15304.n6 a_30192_n15304.n5 10.5449
R18126 a_30192_n15304.n7 a_30192_n15304.n6 10.5449
R18127 a_30192_n15304.n8 a_30192_n15304.n7 10.5449
R18128 a_30192_n15304.n0 a_30192_n15304.t2 10.4819
R18129 a_30192_n15304.n11 a_30192_n15304.n8 8.41578
R18130 a_30192_n15304.n0 a_30192_n15304.n2 7.31398
R18131 a_30192_n15304.n12 a_30192_n15304.n0 6.25311
R18132 a_30192_n15304.n0 a_30192_n15304.n1 5.37659
R18133 a_30192_n15304.n2 a_30192_n15304.t0 4.04494
R18134 a_30192_n15304.n2 a_30192_n15304.t1 4.04494
R18135 a_30192_n15304.n1 a_30192_n15304.t5 3.07367
R18136 a_30192_n15304.n1 a_30192_n15304.t3 3.07367
R18137 a_30192_n15304.n12 a_30192_n15304.t4 3.07367
R18138 a_30192_n15304.t6 a_30192_n15304.n12 3.07367
R18139 a_30192_n15304.n0 a_30192_n15304.n11 2.93567
R18140 a_30192_n15304.n11 a_30192_n15304.n10 2.12967
R18141 a_21772_n17700.n5 a_21772_n17700.t12 15.8415
R18142 a_21772_n17700.n6 a_21772_n17700.t16 15.8415
R18143 a_21772_n17700.n7 a_21772_n17700.t19 15.8415
R18144 a_21772_n17700.n8 a_21772_n17700.t13 15.8415
R18145 a_21772_n17700.n9 a_21772_n17700.t10 15.8415
R18146 a_21772_n17700.n10 a_21772_n17700.t11 15.8415
R18147 a_21772_n17700.n4 a_21772_n17700.t18 15.8415
R18148 a_21772_n17700.n11 a_21772_n17700.t15 15.8415
R18149 a_21772_n17700.n5 a_21772_n17700.t21 13.4447
R18150 a_21772_n17700.n6 a_21772_n17700.t14 13.4447
R18151 a_21772_n17700.n7 a_21772_n17700.t9 13.4447
R18152 a_21772_n17700.n8 a_21772_n17700.t22 13.4447
R18153 a_21772_n17700.n9 a_21772_n17700.t17 13.4447
R18154 a_21772_n17700.n10 a_21772_n17700.t20 13.4447
R18155 a_21772_n17700.n4 a_21772_n17700.t8 13.4447
R18156 a_21772_n17700.n11 a_21772_n17700.t23 13.4447
R18157 a_21772_n17700.n6 a_21772_n17700.n5 10.5449
R18158 a_21772_n17700.n7 a_21772_n17700.n6 10.5449
R18159 a_21772_n17700.n8 a_21772_n17700.n7 10.5449
R18160 a_21772_n17700.n9 a_21772_n17700.n8 10.5449
R18161 a_21772_n17700.n10 a_21772_n17700.n9 10.5449
R18162 a_21772_n17700.n11 a_21772_n17700.n4 10.5449
R18163 a_21772_n17700.n11 a_21772_n17700.n10 10.5449
R18164 a_21772_n17700.n0 a_21772_n17700.n3 7.22489
R18165 a_21772_n17700.n0 a_21772_n17700.n2 6.36702
R18166 a_21772_n17700.n0 a_21772_n17700.n1 3.56115
R18167 a_21772_n17700.n12 a_21772_n17700.n0 2.68463
R18168 a_21772_n17700.n0 a_21772_n17700.n11 2.37183
R18169 a_21772_n17700.n1 a_21772_n17700.t4 2.06607
R18170 a_21772_n17700.n12 a_21772_n17700.t6 2.06607
R18171 a_21772_n17700.n2 a_21772_n17700.t2 1.99806
R18172 a_21772_n17700.n2 a_21772_n17700.t1 1.99806
R18173 a_21772_n17700.n3 a_21772_n17700.t0 1.99806
R18174 a_21772_n17700.n3 a_21772_n17700.t3 1.99806
R18175 a_21772_n17700.n1 a_21772_n17700.t5 1.4923
R18176 a_21772_n17700.t7 a_21772_n17700.n12 1.4923
R18177 a_29744_n15604.n8 a_29744_n15604.t19 15.7685
R18178 a_29744_n15604.n9 a_29744_n15604.t17 15.7685
R18179 a_29744_n15604.n2 a_29744_n15604.t21 15.7685
R18180 a_29744_n15604.n3 a_29744_n15604.t20 15.7685
R18181 a_29744_n15604.n4 a_29744_n15604.t16 15.7685
R18182 a_29744_n15604.n5 a_29744_n15604.t22 15.7685
R18183 a_29744_n15604.n6 a_29744_n15604.t18 15.7685
R18184 a_29744_n15604.n7 a_29744_n15604.t7 15.7685
R18185 a_29744_n15604.n8 a_29744_n15604.t9 11.6197
R18186 a_29744_n15604.n9 a_29744_n15604.t11 11.6197
R18187 a_29744_n15604.n2 a_29744_n15604.t14 11.6197
R18188 a_29744_n15604.n3 a_29744_n15604.t10 11.6197
R18189 a_29744_n15604.n4 a_29744_n15604.t8 11.6197
R18190 a_29744_n15604.n5 a_29744_n15604.t13 11.6197
R18191 a_29744_n15604.n6 a_29744_n15604.t12 11.6197
R18192 a_29744_n15604.n7 a_29744_n15604.t15 11.6197
R18193 a_29744_n15604.n9 a_29744_n15604.n8 10.5449
R18194 a_29744_n15604.n3 a_29744_n15604.n2 10.5449
R18195 a_29744_n15604.n4 a_29744_n15604.n3 10.5449
R18196 a_29744_n15604.n5 a_29744_n15604.n4 10.5449
R18197 a_29744_n15604.n6 a_29744_n15604.n5 10.5449
R18198 a_29744_n15604.n7 a_29744_n15604.n6 10.5449
R18199 a_29744_n15604.n0 a_29744_n15604.t1 10.4819
R18200 a_29744_n15604.n10 a_29744_n15604.n7 8.41578
R18201 a_29744_n15604.n0 a_29744_n15604.n1 7.31398
R18202 a_29744_n15604.n0 a_29744_n15604.n11 6.25311
R18203 a_29744_n15604.n12 a_29744_n15604.n0 5.37659
R18204 a_29744_n15604.n1 a_29744_n15604.t2 4.04494
R18205 a_29744_n15604.n1 a_29744_n15604.t0 4.04494
R18206 a_29744_n15604.n11 a_29744_n15604.t3 3.07367
R18207 a_29744_n15604.n11 a_29744_n15604.t5 3.07367
R18208 a_29744_n15604.n12 a_29744_n15604.t4 3.07367
R18209 a_29744_n15604.t6 a_29744_n15604.n12 3.07367
R18210 a_29744_n15604.n0 a_29744_n15604.n10 2.93567
R18211 a_29744_n15604.n10 a_29744_n15604.n9 2.12967
R18212 a_21772_n14564.n2 a_21772_n14564.t8 15.8415
R18213 a_21772_n14564.n3 a_21772_n14564.t12 15.8415
R18214 a_21772_n14564.n4 a_21772_n14564.t15 15.8415
R18215 a_21772_n14564.n5 a_21772_n14564.t9 15.8415
R18216 a_21772_n14564.n6 a_21772_n14564.t6 15.8415
R18217 a_21772_n14564.n7 a_21772_n14564.t7 15.8415
R18218 a_21772_n14564.n1 a_21772_n14564.t14 15.8415
R18219 a_21772_n14564.n0 a_21772_n14564.t11 15.8415
R18220 a_21772_n14564.n2 a_21772_n14564.t17 13.4447
R18221 a_21772_n14564.n3 a_21772_n14564.t10 13.4447
R18222 a_21772_n14564.n4 a_21772_n14564.t5 13.4447
R18223 a_21772_n14564.n5 a_21772_n14564.t18 13.4447
R18224 a_21772_n14564.n6 a_21772_n14564.t13 13.4447
R18225 a_21772_n14564.n7 a_21772_n14564.t16 13.4447
R18226 a_21772_n14564.n1 a_21772_n14564.t4 13.4447
R18227 a_21772_n14564.n0 a_21772_n14564.t19 13.4447
R18228 a_21772_n14564.n3 a_21772_n14564.n2 10.5449
R18229 a_21772_n14564.n4 a_21772_n14564.n3 10.5449
R18230 a_21772_n14564.n5 a_21772_n14564.n4 10.5449
R18231 a_21772_n14564.n6 a_21772_n14564.n5 10.5449
R18232 a_21772_n14564.n7 a_21772_n14564.n6 10.5449
R18233 a_21772_n14564.n0 a_21772_n14564.n1 10.5449
R18234 a_21772_n14564.n0 a_21772_n14564.n7 10.5449
R18235 a_21772_n14564.n0 a_21772_n14564.t0 7.22489
R18236 a_21772_n14564.t1 a_21772_n14564.n0 7.12153
R18237 a_21772_n14564.n0 a_21772_n14564.t3 6.36702
R18238 a_21772_n14564.n0 a_21772_n14564.t2 5.62673
R18239 a_13623_n12196.n0 a_13623_n12196.t21 56.1018
R18240 a_13623_n12196.n2 a_13623_n12196.t23 56.0719
R18241 a_13623_n12196.n0 a_13623_n12196.t17 56.0141
R18242 a_13623_n12196.n0 a_13623_n12196.t32 55.9719
R18243 a_13623_n12196.n0 a_13623_n12196.t44 55.9719
R18244 a_13623_n12196.n0 a_13623_n12196.t24 55.9719
R18245 a_13623_n12196.n0 a_13623_n12196.t37 55.9719
R18246 a_13623_n12196.n0 a_13623_n12196.t29 55.9719
R18247 a_13623_n12196.n0 a_13623_n12196.t39 55.9719
R18248 a_13623_n12196.n0 a_13623_n12196.t20 55.9719
R18249 a_13623_n12196.n0 a_13623_n12196.t31 55.9719
R18250 a_13623_n12196.n0 a_13623_n12196.t43 55.9719
R18251 a_13623_n12196.n0 a_13623_n12196.t27 55.9719
R18252 a_13623_n12196.n0 a_13623_n12196.t41 55.9719
R18253 a_13623_n12196.n0 a_13623_n12196.t18 55.9719
R18254 a_13623_n12196.n0 a_13623_n12196.t34 55.9719
R18255 a_13623_n12196.n0 a_13623_n12196.t25 55.9719
R18256 a_13623_n12196.n0 a_13623_n12196.t35 55.9719
R18257 a_13623_n12196.n0 a_13623_n12196.t16 55.9719
R18258 a_13623_n12196.n0 a_13623_n12196.t26 55.9719
R18259 a_13623_n12196.n0 a_13623_n12196.t40 55.9719
R18260 a_13623_n12196.n2 a_13623_n12196.t36 55.9719
R18261 a_13623_n12196.n2 a_13623_n12196.t45 55.9719
R18262 a_13623_n12196.n2 a_13623_n12196.t38 55.9719
R18263 a_13623_n12196.n2 a_13623_n12196.t19 55.9719
R18264 a_13623_n12196.n2 a_13623_n12196.t30 55.9719
R18265 a_13623_n12196.n2 a_13623_n12196.t42 55.9719
R18266 a_13623_n12196.n4 a_13623_n12196.t22 55.9719
R18267 a_13623_n12196.n4 a_13623_n12196.t33 55.9719
R18268 a_13623_n12196.n4 a_13623_n12196.t28 55.9719
R18269 a_13623_n12196.n3 a_13623_n12196.n0 32.4358
R18270 a_13623_n12196.n1 a_13623_n12196.n9 6.90733
R18271 a_13623_n12196.n1 a_13623_n12196.n11 6.89497
R18272 a_13623_n12196.n1 a_13623_n12196.n10 6.3768
R18273 a_13623_n12196.n1 a_13623_n12196.n8 6.3768
R18274 a_13623_n12196.n1 a_13623_n12196.n5 3.21104
R18275 a_13623_n12196.n3 a_13623_n12196.n7 2.83209
R18276 a_13623_n12196.n1 a_13623_n12196.n6 2.7042
R18277 a_13623_n12196.n12 a_13623_n12196.n1 2.7042
R18278 a_13623_n12196.n6 a_13623_n12196.t8 2.06607
R18279 a_13623_n12196.n7 a_13623_n12196.t13 2.06607
R18280 a_13623_n12196.n5 a_13623_n12196.t9 2.06607
R18281 a_13623_n12196.t15 a_13623_n12196.n12 2.06607
R18282 a_13623_n12196.n10 a_13623_n12196.t3 1.99806
R18283 a_13623_n12196.n10 a_13623_n12196.t4 1.99806
R18284 a_13623_n12196.n11 a_13623_n12196.t7 1.99806
R18285 a_13623_n12196.n11 a_13623_n12196.t0 1.99806
R18286 a_13623_n12196.n9 a_13623_n12196.t5 1.99806
R18287 a_13623_n12196.n9 a_13623_n12196.t2 1.99806
R18288 a_13623_n12196.n8 a_13623_n12196.t1 1.99806
R18289 a_13623_n12196.n8 a_13623_n12196.t6 1.99806
R18290 a_13623_n12196.n6 a_13623_n12196.t12 1.4923
R18291 a_13623_n12196.n7 a_13623_n12196.t10 1.4923
R18292 a_13623_n12196.n5 a_13623_n12196.t11 1.4923
R18293 a_13623_n12196.n12 a_13623_n12196.t14 1.4923
R18294 a_13623_n12196.n1 a_13623_n12196.n3 1.23036
R18295 a_13623_n12196.n0 a_13623_n12196.n4 1.21355
R18296 a_13623_n12196.n4 a_13623_n12196.n2 0.8005
R18297 CLK CLK.n7 40.9248
R18298 CLK.n1 CLK.t15 31.7717
R18299 CLK.n3 CLK.t4 29.7439
R18300 CLK.n3 CLK.t2 18.7615
R18301 CLK.n4 CLK.t5 18.7615
R18302 CLK.n5 CLK.t11 18.7615
R18303 CLK.n1 CLK.t8 18.7615
R18304 CLK.n2 CLK.t9 18.7615
R18305 CLK.n6 CLK.t7 18.7615
R18306 CLK.n3 CLK.t10 11.133
R18307 CLK.n4 CLK.t13 11.133
R18308 CLK.n5 CLK.t14 11.133
R18309 CLK.n1 CLK.t1 11.133
R18310 CLK.n2 CLK.t3 11.133
R18311 CLK.n6 CLK.t0 11.133
R18312 CLK.n4 CLK.n3 10.5449
R18313 CLK.n5 CLK.n4 10.5449
R18314 CLK.n2 CLK.n1 10.5449
R18315 CLK.n6 CLK.n2 10.5449
R18316 CLK.n6 CLK.n5 10.5449
R18317 CLK.n0 CLK.t6 6.56378
R18318 CLK.n7 CLK.n6 6.50965
R18319 CLK.n0 CLK.t12 5.35632
R18320 CLK.n7 CLK.n0 4.5005
R18321 a_24348_n16087.n2 a_24348_n16087.n0 31.7018
R18322 a_24348_n16087.n1 a_24348_n16087.t5 29.2005
R18323 a_24348_n16087.n3 a_24348_n16087.t3 19.7105
R18324 a_24348_n16087.n0 a_24348_n16087.t2 19.0535
R18325 a_24348_n16087.n4 a_24348_n16087.n3 17.4744
R18326 a_24348_n16087.n2 a_24348_n16087.n1 13.7886
R18327 a_24348_n16087.n3 a_24348_n16087.t6 13.3108
R18328 a_24348_n16087.n1 a_24348_n16087.t7 12.1428
R18329 a_24348_n16087.n0 a_24348_n16087.t4 10.9505
R18330 a_24348_n16087.t1 a_24348_n16087.n4 9.02222
R18331 a_24348_n16087.t1 a_24348_n16087.t0 8.76859
R18332 a_24348_n16087.n4 a_24348_n16087.n2 7.0205
R18333 a_13623_n14874.n0 a_13623_n14874.t43 56.1018
R18334 a_13623_n14874.n2 a_13623_n14874.t22 56.0719
R18335 a_13623_n14874.n0 a_13623_n14874.t17 56.0141
R18336 a_13623_n14874.n0 a_13623_n14874.t24 55.9719
R18337 a_13623_n14874.n0 a_13623_n14874.t37 55.9719
R18338 a_13623_n14874.n0 a_13623_n14874.t45 55.9719
R18339 a_13623_n14874.n0 a_13623_n14874.t29 55.9719
R18340 a_13623_n14874.n0 a_13623_n14874.t20 55.9719
R18341 a_13623_n14874.n0 a_13623_n14874.t31 55.9719
R18342 a_13623_n14874.n0 a_13623_n14874.t42 55.9719
R18343 a_13623_n14874.n0 a_13623_n14874.t23 55.9719
R18344 a_13623_n14874.n0 a_13623_n14874.t36 55.9719
R18345 a_13623_n14874.n0 a_13623_n14874.t27 55.9719
R18346 a_13623_n14874.n0 a_13623_n14874.t40 55.9719
R18347 a_13623_n14874.n0 a_13623_n14874.t18 55.9719
R18348 a_13623_n14874.n0 a_13623_n14874.t33 55.9719
R18349 a_13623_n14874.n0 a_13623_n14874.t25 55.9719
R18350 a_13623_n14874.n0 a_13623_n14874.t34 55.9719
R18351 a_13623_n14874.n0 a_13623_n14874.t16 55.9719
R18352 a_13623_n14874.n0 a_13623_n14874.t26 55.9719
R18353 a_13623_n14874.n0 a_13623_n14874.t39 55.9719
R18354 a_13623_n14874.n2 a_13623_n14874.t35 55.9719
R18355 a_13623_n14874.n2 a_13623_n14874.t44 55.9719
R18356 a_13623_n14874.n2 a_13623_n14874.t38 55.9719
R18357 a_13623_n14874.n2 a_13623_n14874.t19 55.9719
R18358 a_13623_n14874.n2 a_13623_n14874.t30 55.9719
R18359 a_13623_n14874.n2 a_13623_n14874.t41 55.9719
R18360 a_13623_n14874.n4 a_13623_n14874.t21 55.9719
R18361 a_13623_n14874.n4 a_13623_n14874.t32 55.9719
R18362 a_13623_n14874.n4 a_13623_n14874.t28 55.9719
R18363 a_13623_n14874.n3 a_13623_n14874.n0 32.2815
R18364 a_13623_n14874.n1 a_13623_n14874.n9 6.90733
R18365 a_13623_n14874.n1 a_13623_n14874.n11 6.89497
R18366 a_13623_n14874.n1 a_13623_n14874.n10 6.3768
R18367 a_13623_n14874.n1 a_13623_n14874.n8 6.3768
R18368 a_13623_n14874.n1 a_13623_n14874.n5 3.21104
R18369 a_13623_n14874.n3 a_13623_n14874.n7 2.83209
R18370 a_13623_n14874.n1 a_13623_n14874.n6 2.7042
R18371 a_13623_n14874.n12 a_13623_n14874.n1 2.7042
R18372 a_13623_n14874.n6 a_13623_n14874.t8 2.06607
R18373 a_13623_n14874.n7 a_13623_n14874.t13 2.06607
R18374 a_13623_n14874.n5 a_13623_n14874.t9 2.06607
R18375 a_13623_n14874.t15 a_13623_n14874.n12 2.06607
R18376 a_13623_n14874.n10 a_13623_n14874.t5 1.99806
R18377 a_13623_n14874.n10 a_13623_n14874.t6 1.99806
R18378 a_13623_n14874.n11 a_13623_n14874.t1 1.99806
R18379 a_13623_n14874.n11 a_13623_n14874.t2 1.99806
R18380 a_13623_n14874.n9 a_13623_n14874.t7 1.99806
R18381 a_13623_n14874.n9 a_13623_n14874.t4 1.99806
R18382 a_13623_n14874.n8 a_13623_n14874.t3 1.99806
R18383 a_13623_n14874.n8 a_13623_n14874.t0 1.99806
R18384 a_13623_n14874.n6 a_13623_n14874.t12 1.4923
R18385 a_13623_n14874.n7 a_13623_n14874.t10 1.4923
R18386 a_13623_n14874.n5 a_13623_n14874.t11 1.4923
R18387 a_13623_n14874.n12 a_13623_n14874.t14 1.4923
R18388 a_13623_n14874.n1 a_13623_n14874.n3 1.23036
R18389 a_13623_n14874.n0 a_13623_n14874.n4 1.21355
R18390 a_13623_n14874.n4 a_13623_n14874.n2 0.8005
R18391 a_37024_1944.n10 a_37024_1944.t8 15.8415
R18392 a_37024_1944.n4 a_37024_1944.t11 15.8415
R18393 a_37024_1944.n5 a_37024_1944.t14 15.8415
R18394 a_37024_1944.n6 a_37024_1944.t9 15.8415
R18395 a_37024_1944.n7 a_37024_1944.t23 15.8415
R18396 a_37024_1944.n8 a_37024_1944.t13 15.8415
R18397 a_37024_1944.n9 a_37024_1944.t10 15.8415
R18398 a_37024_1944.n11 a_37024_1944.t12 15.8415
R18399 a_37024_1944.n10 a_37024_1944.t16 13.4447
R18400 a_37024_1944.n4 a_37024_1944.t19 13.4447
R18401 a_37024_1944.n5 a_37024_1944.t22 13.4447
R18402 a_37024_1944.n6 a_37024_1944.t17 13.4447
R18403 a_37024_1944.n7 a_37024_1944.t15 13.4447
R18404 a_37024_1944.n8 a_37024_1944.t21 13.4447
R18405 a_37024_1944.n9 a_37024_1944.t18 13.4447
R18406 a_37024_1944.n11 a_37024_1944.t20 13.4447
R18407 a_37024_1944.n5 a_37024_1944.n4 10.5449
R18408 a_37024_1944.n6 a_37024_1944.n5 10.5449
R18409 a_37024_1944.n7 a_37024_1944.n6 10.5449
R18410 a_37024_1944.n8 a_37024_1944.n7 10.5449
R18411 a_37024_1944.n9 a_37024_1944.n8 10.5449
R18412 a_37024_1944.n11 a_37024_1944.n9 10.5449
R18413 a_37024_1944.n11 a_37024_1944.n10 10.5449
R18414 a_37024_1944.n0 a_37024_1944.n3 7.22489
R18415 a_37024_1944.n0 a_37024_1944.n2 6.36702
R18416 a_37024_1944.n12 a_37024_1944.n0 3.56115
R18417 a_37024_1944.n0 a_37024_1944.n1 2.68463
R18418 a_37024_1944.n0 a_37024_1944.n11 2.37181
R18419 a_37024_1944.n1 a_37024_1944.t6 2.06607
R18420 a_37024_1944.t7 a_37024_1944.n12 2.06607
R18421 a_37024_1944.n2 a_37024_1944.t1 1.99806
R18422 a_37024_1944.n2 a_37024_1944.t0 1.99806
R18423 a_37024_1944.n3 a_37024_1944.t2 1.99806
R18424 a_37024_1944.n3 a_37024_1944.t3 1.99806
R18425 a_37024_1944.n1 a_37024_1944.t5 1.4923
R18426 a_37024_1944.n12 a_37024_1944.t4 1.4923
R18427 OUT[2] OUT[2].n14 22.8425
R18428 OUT[2].n3 OUT[2].n2 6.90733
R18429 OUT[2].n3 OUT[2].n1 6.3768
R18430 OUT[2].n12 OUT[2].n0 6.3768
R18431 OUT[2].n14 OUT[2].n13 6.3005
R18432 OUT[2].n9 OUT[2].n8 3.23472
R18433 OUT[2].n6 OUT[2].n5 3.21104
R18434 OUT[2].n9 OUT[2].n7 2.7042
R18435 OUT[2].n6 OUT[2].n4 2.7042
R18436 OUT[2].n7 OUT[2].t14 2.06607
R18437 OUT[2].n8 OUT[2].t12 2.06607
R18438 OUT[2].n5 OUT[2].t15 2.06607
R18439 OUT[2].n4 OUT[2].t10 2.06607
R18440 OUT[2].n13 OUT[2].t2 1.99806
R18441 OUT[2].n13 OUT[2].t6 1.99806
R18442 OUT[2].n2 OUT[2].t3 1.99806
R18443 OUT[2].n2 OUT[2].t0 1.99806
R18444 OUT[2].n1 OUT[2].t5 1.99806
R18445 OUT[2].n1 OUT[2].t7 1.99806
R18446 OUT[2].n0 OUT[2].t1 1.99806
R18447 OUT[2].n0 OUT[2].t4 1.99806
R18448 OUT[2].n7 OUT[2].t8 1.4923
R18449 OUT[2].n8 OUT[2].t9 1.4923
R18450 OUT[2].n5 OUT[2].t11 1.4923
R18451 OUT[2].n4 OUT[2].t13 1.4923
R18452 OUT[2].n14 OUT[2].n12 0.577837
R18453 OUT[2].n11 OUT[2].n3 0.189974
R18454 OUT[2].n10 OUT[2].n6 0.175763
R18455 OUT[2].n10 OUT[2].n9 0.166289
R18456 OUT[2].n12 OUT[2].n11 0.152079
R18457 OUT[2].n11 OUT[2].n10 0.145625
R18458 a_11023_n20230.n21 a_11023_n20230.t30 56.0276
R18459 a_11023_n20230.n10 a_11023_n20230.t32 56.019
R18460 a_11023_n20230.n12 a_11023_n20230.t28 55.9719
R18461 a_11023_n20230.n6 a_11023_n20230.t36 55.9719
R18462 a_11023_n20230.n14 a_11023_n20230.t23 55.9719
R18463 a_11023_n20230.n5 a_11023_n20230.t38 55.9719
R18464 a_11023_n20230.n16 a_11023_n20230.t24 55.9719
R18465 a_11023_n20230.n4 a_11023_n20230.t33 55.9719
R18466 a_11023_n20230.n17 a_11023_n20230.t21 55.9719
R18467 a_11023_n20230.n2 a_11023_n20230.t27 55.9719
R18468 a_11023_n20230.n22 a_11023_n20230.t35 55.9719
R18469 a_11023_n20230.n10 a_11023_n20230.t20 55.9719
R18470 a_11023_n20230.n10 a_11023_n20230.t26 55.9719
R18471 a_11023_n20230.n9 a_11023_n20230.t34 55.9719
R18472 a_11023_n20230.n9 a_11023_n20230.t22 55.9719
R18473 a_11023_n20230.n7 a_11023_n20230.t29 55.9719
R18474 a_11023_n20230.n7 a_11023_n20230.t37 55.9719
R18475 a_11023_n20230.n8 a_11023_n20230.t31 55.9719
R18476 a_11023_n20230.n8 a_11023_n20230.t39 55.9719
R18477 a_11023_n20230.n27 a_11023_n20230.t25 55.9719
R18478 a_11023_n20230.n12 a_11023_n20230.n11 0.0590857
R18479 a_11023_n20230.n24 a_11023_n20230.n23 4.5005
R18480 a_11023_n20230.n25 a_11023_n20230.n2 4.5005
R18481 a_11023_n20230.n17 a_11023_n20230.n26 4.5005
R18482 a_11023_n20230.n3 a_11023_n20230.n0 4.5005
R18483 a_11023_n20230.n1 a_11023_n20230.n4 4.5005
R18484 a_11023_n20230.n16 a_11023_n20230.n15 4.5005
R18485 a_11023_n20230.n33 a_11023_n20230.n32 4.5005
R18486 a_11023_n20230.n31 a_11023_n20230.n5 4.5005
R18487 a_11023_n20230.n14 a_11023_n20230.n13 4.5005
R18488 a_11023_n20230.n30 a_11023_n20230.n29 4.5005
R18489 a_11023_n20230.n28 a_11023_n20230.n6 4.5005
R18490 a_11023_n20230.n39 a_11023_n20230.n38 3.87048
R18491 a_11023_n20230.n39 a_11023_n20230.n37 3.68704
R18492 a_11023_n20230.n40 a_11023_n20230.n36 3.68704
R18493 a_11023_n20230.n41 a_11023_n20230.n35 3.68704
R18494 a_11023_n20230.n42 a_11023_n20230.n34 3.68704
R18495 a_11023_n20230.n20 a_11023_n20230.n18 3.53719
R18496 a_11023_n20230.n45 a_11023_n20230.n44 3.37808
R18497 a_11023_n20230.n47 a_11023_n20230.n46 3.37808
R18498 a_11023_n20230.n20 a_11023_n20230.n19 3.37808
R18499 a_11023_n20230.n49 a_11023_n20230.n48 3.37783
R18500 a_11023_n20230.n43 a_11023_n20230.n1 1.89107
R18501 a_11023_n20230.n24 a_11023_n20230.n21 1.15666
R18502 a_11023_n20230.n44 a_11023_n20230.t10 0.6505
R18503 a_11023_n20230.n44 a_11023_n20230.t14 0.6505
R18504 a_11023_n20230.n46 a_11023_n20230.t13 0.6505
R18505 a_11023_n20230.n46 a_11023_n20230.t16 0.6505
R18506 a_11023_n20230.n19 a_11023_n20230.t15 0.6505
R18507 a_11023_n20230.n19 a_11023_n20230.t18 0.6505
R18508 a_11023_n20230.n18 a_11023_n20230.t17 0.6505
R18509 a_11023_n20230.n18 a_11023_n20230.t11 0.6505
R18510 a_11023_n20230.n49 a_11023_n20230.t12 0.6505
R18511 a_11023_n20230.t19 a_11023_n20230.n49 0.6505
R18512 a_11023_n20230.n38 a_11023_n20230.t5 0.5855
R18513 a_11023_n20230.n38 a_11023_n20230.t9 0.5855
R18514 a_11023_n20230.n37 a_11023_n20230.t3 0.5855
R18515 a_11023_n20230.n37 a_11023_n20230.t6 0.5855
R18516 a_11023_n20230.n36 a_11023_n20230.t0 0.5855
R18517 a_11023_n20230.n36 a_11023_n20230.t7 0.5855
R18518 a_11023_n20230.n35 a_11023_n20230.t1 0.5855
R18519 a_11023_n20230.n35 a_11023_n20230.t4 0.5855
R18520 a_11023_n20230.n34 a_11023_n20230.t8 0.5855
R18521 a_11023_n20230.n34 a_11023_n20230.t2 0.5855
R18522 a_11023_n20230.n43 a_11023_n20230.n42 0.41138
R18523 a_11023_n20230.n45 a_11023_n20230.n43 0.373278
R18524 a_11023_n20230.n40 a_11023_n20230.n39 0.183939
R18525 a_11023_n20230.n41 a_11023_n20230.n40 0.183939
R18526 a_11023_n20230.n42 a_11023_n20230.n41 0.183939
R18527 a_11023_n20230.n48 a_11023_n20230.n20 0.159616
R18528 a_11023_n20230.n48 a_11023_n20230.n47 0.159616
R18529 a_11023_n20230.n47 a_11023_n20230.n45 0.159616
R18530 a_11023_n20230.n22 a_11023_n20230.n21 0.121859
R18531 a_11023_n20230.n23 a_11023_n20230.n22 0.11975
R18532 a_11023_n20230.n17 a_11023_n20230.n2 0.11975
R18533 a_11023_n20230.n4 a_11023_n20230.n16 0.11975
R18534 a_11023_n20230.n5 a_11023_n20230.n14 0.11975
R18535 a_11023_n20230.n6 a_11023_n20230.n12 0.11975
R18536 a_11023_n20230.n25 a_11023_n20230.n24 0.11975
R18537 a_11023_n20230.n26 a_11023_n20230.n25 0.11975
R18538 a_11023_n20230.n26 a_11023_n20230.n0 0.11975
R18539 a_11023_n20230.n1 a_11023_n20230.n15 0.11975
R18540 a_11023_n20230.n32 a_11023_n20230.n15 0.11975
R18541 a_11023_n20230.n32 a_11023_n20230.n31 0.11975
R18542 a_11023_n20230.n31 a_11023_n20230.n13 0.11975
R18543 a_11023_n20230.n29 a_11023_n20230.n13 0.11975
R18544 a_11023_n20230.n29 a_11023_n20230.n28 0.11975
R18545 a_11023_n20230.n28 a_11023_n20230.n11 2.37025
R18546 a_11023_n20230.n3 a_11023_n20230.n17 0.11975
R18547 a_11023_n20230.n16 a_11023_n20230.n33 0.11975
R18548 a_11023_n20230.n14 a_11023_n20230.n30 0.11975
R18549 a_11023_n20230.n11 a_11023_n20230.n27 1.35571
R18550 a_11023_n20230.n30 a_11023_n20230.n6 0.11975
R18551 a_11023_n20230.n33 a_11023_n20230.n5 0.11975
R18552 a_11023_n20230.n4 a_11023_n20230.n3 0.11975
R18553 a_11023_n20230.n23 a_11023_n20230.n2 0.11975
R18554 a_11023_n20230.n1 a_11023_n20230.n0 0.11975
R18555 a_11023_n20230.n9 a_11023_n20230.n10 0.0946176
R18556 a_11023_n20230.n7 a_11023_n20230.n9 0.0946176
R18557 a_11023_n20230.n8 a_11023_n20230.n7 0.0946176
R18558 a_11023_n20230.n27 a_11023_n20230.n8 0.0946176
R18559 a_1955_4292.n0 a_1955_4292.t2 61.8885
R18560 a_1955_4292.n0 a_1955_4292.t4 60.7348
R18561 a_1955_4292.n1 a_1955_4292.t3 56.2348
R18562 a_1955_4292.n2 a_1955_4292.n1 16.4203
R18563 a_1955_4292.n1 a_1955_4292.n0 5.4365
R18564 a_1955_4292.n2 a_1955_4292.t1 2.96547
R18565 a_1955_4292.t0 a_1955_4292.n2 2.5601
R18566 a_24236_2258.t1 a_24236_2258.n3 53.2582
R18567 a_24236_2258.n2 a_24236_2258.t5 17.119
R18568 a_24236_2258.n0 a_24236_2258.t8 16.2065
R18569 a_24236_2258.n1 a_24236_2258.t2 16.2065
R18570 a_24236_2258.n3 a_24236_2258.t4 16.2065
R18571 a_24236_2258.n1 a_24236_2258.t3 13.1405
R18572 a_24236_2258.n3 a_24236_2258.t7 13.1405
R18573 a_24236_2258.n2 a_24236_2258.t6 12.228
R18574 a_24236_2258.n0 a_24236_2258.t9 12.228
R18575 a_24236_2258.n3 a_24236_2258.n1 10.5449
R18576 a_24236_2258.n3 a_24236_2258.n0 10.5449
R18577 a_24236_2258.t1 a_24236_2258.t0 9.70112
R18578 a_24236_2258.n0 a_24236_2258.n2 8.35614
R18579 a_22444_2253.n5 a_22444_2253.t11 15.8415
R18580 a_22444_2253.n6 a_22444_2253.t9 15.8415
R18581 a_22444_2253.n7 a_22444_2253.t8 15.8415
R18582 a_22444_2253.n8 a_22444_2253.t13 15.8415
R18583 a_22444_2253.n9 a_22444_2253.t19 15.8415
R18584 a_22444_2253.n10 a_22444_2253.t15 15.8415
R18585 a_22444_2253.n4 a_22444_2253.t20 15.8415
R18586 a_22444_2253.n11 a_22444_2253.t23 15.8415
R18587 a_22444_2253.n5 a_22444_2253.t14 13.4447
R18588 a_22444_2253.n6 a_22444_2253.t10 13.4447
R18589 a_22444_2253.n7 a_22444_2253.t17 13.4447
R18590 a_22444_2253.n8 a_22444_2253.t16 13.4447
R18591 a_22444_2253.n9 a_22444_2253.t21 13.4447
R18592 a_22444_2253.n10 a_22444_2253.t18 13.4447
R18593 a_22444_2253.n4 a_22444_2253.t22 13.4447
R18594 a_22444_2253.n11 a_22444_2253.t12 13.4447
R18595 a_22444_2253.n6 a_22444_2253.n5 10.5449
R18596 a_22444_2253.n7 a_22444_2253.n6 10.5449
R18597 a_22444_2253.n8 a_22444_2253.n7 10.5449
R18598 a_22444_2253.n9 a_22444_2253.n8 10.5449
R18599 a_22444_2253.n10 a_22444_2253.n9 10.5449
R18600 a_22444_2253.n11 a_22444_2253.n4 10.5449
R18601 a_22444_2253.n11 a_22444_2253.n10 10.5449
R18602 a_22444_2253.n0 a_22444_2253.n3 7.22489
R18603 a_22444_2253.n0 a_22444_2253.n2 6.36702
R18604 a_22444_2253.n12 a_22444_2253.n0 3.56115
R18605 a_22444_2253.n0 a_22444_2253.n1 2.68463
R18606 a_22444_2253.n0 a_22444_2253.n11 2.37048
R18607 a_22444_2253.n1 a_22444_2253.t5 2.06607
R18608 a_22444_2253.n12 a_22444_2253.t6 2.06607
R18609 a_22444_2253.n3 a_22444_2253.t3 1.99806
R18610 a_22444_2253.n3 a_22444_2253.t1 1.99806
R18611 a_22444_2253.n2 a_22444_2253.t0 1.99806
R18612 a_22444_2253.n2 a_22444_2253.t2 1.99806
R18613 a_22444_2253.n1 a_22444_2253.t4 1.4923
R18614 a_22444_2253.t7 a_22444_2253.n12 1.4923
R18615 a_29408_1944.n10 a_29408_1944.t19 15.8415
R18616 a_29408_1944.n4 a_29408_1944.t22 15.8415
R18617 a_29408_1944.n5 a_29408_1944.t18 15.8415
R18618 a_29408_1944.n6 a_29408_1944.t21 15.8415
R18619 a_29408_1944.n7 a_29408_1944.t23 15.8415
R18620 a_29408_1944.n8 a_29408_1944.t17 15.8415
R18621 a_29408_1944.n9 a_29408_1944.t20 15.8415
R18622 a_29408_1944.n11 a_29408_1944.t16 15.8415
R18623 a_29408_1944.n10 a_29408_1944.t11 13.4447
R18624 a_29408_1944.n4 a_29408_1944.t14 13.4447
R18625 a_29408_1944.n5 a_29408_1944.t10 13.4447
R18626 a_29408_1944.n6 a_29408_1944.t13 13.4447
R18627 a_29408_1944.n7 a_29408_1944.t15 13.4447
R18628 a_29408_1944.n8 a_29408_1944.t9 13.4447
R18629 a_29408_1944.n9 a_29408_1944.t12 13.4447
R18630 a_29408_1944.n11 a_29408_1944.t8 13.4447
R18631 a_29408_1944.n5 a_29408_1944.n4 10.5449
R18632 a_29408_1944.n6 a_29408_1944.n5 10.5449
R18633 a_29408_1944.n7 a_29408_1944.n6 10.5449
R18634 a_29408_1944.n8 a_29408_1944.n7 10.5449
R18635 a_29408_1944.n9 a_29408_1944.n8 10.5449
R18636 a_29408_1944.n11 a_29408_1944.n9 10.5449
R18637 a_29408_1944.n11 a_29408_1944.n10 10.5449
R18638 a_29408_1944.n0 a_29408_1944.n3 7.22489
R18639 a_29408_1944.n0 a_29408_1944.n2 6.36702
R18640 a_29408_1944.n12 a_29408_1944.n0 3.56115
R18641 a_29408_1944.n0 a_29408_1944.n1 2.68463
R18642 a_29408_1944.n0 a_29408_1944.n11 2.37181
R18643 a_29408_1944.n1 a_29408_1944.t4 2.06607
R18644 a_29408_1944.n12 a_29408_1944.t5 2.06607
R18645 a_29408_1944.n2 a_29408_1944.t0 1.99806
R18646 a_29408_1944.n2 a_29408_1944.t2 1.99806
R18647 a_29408_1944.n3 a_29408_1944.t1 1.99806
R18648 a_29408_1944.n3 a_29408_1944.t3 1.99806
R18649 a_29408_1944.n1 a_29408_1944.t6 1.4923
R18650 a_29408_1944.t7 a_29408_1944.n12 1.4923
R18651 OUT[0] OUT[0].n14 20.4125
R18652 OUT[0].n3 OUT[0].n2 6.90733
R18653 OUT[0].n3 OUT[0].n1 6.3768
R18654 OUT[0].n12 OUT[0].n0 6.3768
R18655 OUT[0].n14 OUT[0].n13 6.3005
R18656 OUT[0].n9 OUT[0].n8 3.23472
R18657 OUT[0].n6 OUT[0].n5 3.21104
R18658 OUT[0].n9 OUT[0].n7 2.7042
R18659 OUT[0].n6 OUT[0].n4 2.7042
R18660 OUT[0].n7 OUT[0].t10 2.06607
R18661 OUT[0].n8 OUT[0].t9 2.06607
R18662 OUT[0].n5 OUT[0].t12 2.06607
R18663 OUT[0].n4 OUT[0].t14 2.06607
R18664 OUT[0].n13 OUT[0].t7 1.99806
R18665 OUT[0].n13 OUT[0].t4 1.99806
R18666 OUT[0].n2 OUT[0].t1 1.99806
R18667 OUT[0].n2 OUT[0].t5 1.99806
R18668 OUT[0].n1 OUT[0].t2 1.99806
R18669 OUT[0].n1 OUT[0].t0 1.99806
R18670 OUT[0].n0 OUT[0].t6 1.99806
R18671 OUT[0].n0 OUT[0].t3 1.99806
R18672 OUT[0].n7 OUT[0].t8 1.4923
R18673 OUT[0].n8 OUT[0].t13 1.4923
R18674 OUT[0].n5 OUT[0].t15 1.4923
R18675 OUT[0].n4 OUT[0].t11 1.4923
R18676 OUT[0].n14 OUT[0].n12 0.577837
R18677 OUT[0].n11 OUT[0].n3 0.189974
R18678 OUT[0].n10 OUT[0].n6 0.175763
R18679 OUT[0].n10 OUT[0].n9 0.166289
R18680 OUT[0].n12 OUT[0].n11 0.152079
R18681 OUT[0].n11 OUT[0].n10 0.145625
R18682 a_29532_n4372.n5 a_29532_n4372.n1 36.5505
R18683 a_29532_n4372.n3 a_29532_n4372.t6 23.5552
R18684 a_29532_n4372.n2 a_29532_n4372.t9 17.4475
R18685 a_29532_n4372.n2 a_29532_n4372.t8 16.4012
R18686 a_29532_n4372.n1 a_29532_n4372.t5 15.9023
R18687 a_29532_n4372.n1 a_29532_n4372.t7 13.4447
R18688 a_29532_n4372.n0 a_29532_n4372.n5 11.8805
R18689 a_29532_n4372.n3 a_29532_n4372.t4 10.2935
R18690 a_29532_n4372.n4 a_29532_n4372.n3 10.2927
R18691 a_29532_n4372.n4 a_29532_n4372.n2 8.20326
R18692 a_29532_n4372.n0 a_29532_n4372.t2 7.22707
R18693 a_29532_n4372.n0 a_29532_n4372.t3 6.9805
R18694 a_29532_n4372.n0 a_29532_n4372.t0 5.98178
R18695 a_29532_n4372.t1 a_29532_n4372.n0 5.2005
R18696 a_29532_n4372.n5 a_29532_n4372.n4 4.5005
R18697 a_41392_1944.n10 a_41392_1944.t14 15.8415
R18698 a_41392_1944.n4 a_41392_1944.t10 15.8415
R18699 a_41392_1944.n5 a_41392_1944.t13 15.8415
R18700 a_41392_1944.n6 a_41392_1944.t9 15.8415
R18701 a_41392_1944.n7 a_41392_1944.t15 15.8415
R18702 a_41392_1944.n8 a_41392_1944.t12 15.8415
R18703 a_41392_1944.n9 a_41392_1944.t8 15.8415
R18704 a_41392_1944.n11 a_41392_1944.t11 15.8415
R18705 a_41392_1944.n10 a_41392_1944.t22 13.4447
R18706 a_41392_1944.n4 a_41392_1944.t18 13.4447
R18707 a_41392_1944.n5 a_41392_1944.t21 13.4447
R18708 a_41392_1944.n6 a_41392_1944.t17 13.4447
R18709 a_41392_1944.n7 a_41392_1944.t23 13.4447
R18710 a_41392_1944.n8 a_41392_1944.t20 13.4447
R18711 a_41392_1944.n9 a_41392_1944.t16 13.4447
R18712 a_41392_1944.n11 a_41392_1944.t19 13.4447
R18713 a_41392_1944.n5 a_41392_1944.n4 10.5449
R18714 a_41392_1944.n6 a_41392_1944.n5 10.5449
R18715 a_41392_1944.n7 a_41392_1944.n6 10.5449
R18716 a_41392_1944.n8 a_41392_1944.n7 10.5449
R18717 a_41392_1944.n9 a_41392_1944.n8 10.5449
R18718 a_41392_1944.n11 a_41392_1944.n9 10.5449
R18719 a_41392_1944.n11 a_41392_1944.n10 10.5449
R18720 a_41392_1944.n0 a_41392_1944.n3 7.22489
R18721 a_41392_1944.n0 a_41392_1944.n2 6.36702
R18722 a_41392_1944.n12 a_41392_1944.n0 3.56115
R18723 a_41392_1944.n0 a_41392_1944.n1 2.68463
R18724 a_41392_1944.n0 a_41392_1944.n11 2.37181
R18725 a_41392_1944.n1 a_41392_1944.t6 2.06607
R18726 a_41392_1944.t7 a_41392_1944.n12 2.06607
R18727 a_41392_1944.n2 a_41392_1944.t2 1.99806
R18728 a_41392_1944.n2 a_41392_1944.t1 1.99806
R18729 a_41392_1944.n3 a_41392_1944.t3 1.99806
R18730 a_41392_1944.n3 a_41392_1944.t0 1.99806
R18731 a_41392_1944.n1 a_41392_1944.t5 1.4923
R18732 a_41392_1944.n12 a_41392_1944.t4 1.4923
R18733 a_13501_n19850.n1 a_13501_n19850.t10 15.8618
R18734 a_13501_n19850.n0 a_13501_n19850.t19 15.8393
R18735 a_13501_n19850.n1 a_13501_n19850.t5 15.7537
R18736 a_13501_n19850.n0 a_13501_n19850.t4 15.7496
R18737 a_13501_n19850.n0 a_13501_n19850.n2 14.963
R18738 a_13501_n19850.n1 a_13501_n19850.n4 14.9583
R18739 a_13501_n19850.n1 a_13501_n19850.n6 14.9559
R18740 a_13501_n19850.n1 a_13501_n19850.n7 14.9547
R18741 a_13501_n19850.n0 a_13501_n19850.n3 14.7096
R18742 a_13501_n19850.n9 a_13501_n19850.n1 14.7035
R18743 a_13501_n19850.n1 a_13501_n19850.n8 14.7035
R18744 a_13501_n19850.n1 a_13501_n19850.n5 14.6941
R18745 a_13501_n19850.n5 a_13501_n19850.t8 0.6505
R18746 a_13501_n19850.n5 a_13501_n19850.t1 0.6505
R18747 a_13501_n19850.n8 a_13501_n19850.t7 0.6505
R18748 a_13501_n19850.n8 a_13501_n19850.t0 0.6505
R18749 a_13501_n19850.n3 a_13501_n19850.t2 0.6505
R18750 a_13501_n19850.n3 a_13501_n19850.t6 0.6505
R18751 a_13501_n19850.t9 a_13501_n19850.n9 0.6505
R18752 a_13501_n19850.n9 a_13501_n19850.t3 0.6505
R18753 a_13501_n19850.n6 a_13501_n19850.t13 0.5855
R18754 a_13501_n19850.n6 a_13501_n19850.t16 0.5855
R18755 a_13501_n19850.n7 a_13501_n19850.t12 0.5855
R18756 a_13501_n19850.n7 a_13501_n19850.t15 0.5855
R18757 a_13501_n19850.n4 a_13501_n19850.t14 0.5855
R18758 a_13501_n19850.n4 a_13501_n19850.t18 0.5855
R18759 a_13501_n19850.n2 a_13501_n19850.t17 0.5855
R18760 a_13501_n19850.n2 a_13501_n19850.t11 0.5855
R18761 a_13501_n19850.n1 a_13501_n19850.n0 0.158862
R18762 a_n263_3472.n10 a_n263_3472.t16 60.8271
R18763 a_n263_3472.n9 a_n263_3472.t17 56.8971
R18764 a_n263_3472.n9 a_n263_3472.t18 56.5155
R18765 a_n263_3472.n0 a_n263_3472.n10 39.4859
R18766 a_n263_3472.n0 a_n263_3472.n5 6.90733
R18767 a_n263_3472.n1 a_n263_3472.n7 6.89497
R18768 a_n263_3472.n1 a_n263_3472.n6 6.3768
R18769 a_n263_3472.n0 a_n263_3472.n4 6.3768
R18770 a_n263_3472.n10 a_n263_3472.n9 5.5475
R18771 a_n263_3472.n0 a_n263_3472.n3 3.21104
R18772 a_n263_3472.n0 a_n263_3472.n2 2.7042
R18773 a_n263_3472.n0 a_n263_3472.n8 2.7042
R18774 a_n263_3472.n11 a_n263_3472.n0 2.7042
R18775 a_n263_3472.n2 a_n263_3472.t10 2.06607
R18776 a_n263_3472.n3 a_n263_3472.t9 2.06607
R18777 a_n263_3472.n8 a_n263_3472.t13 2.06607
R18778 a_n263_3472.t15 a_n263_3472.n11 2.06607
R18779 a_n263_3472.n7 a_n263_3472.t0 1.99806
R18780 a_n263_3472.n7 a_n263_3472.t6 1.99806
R18781 a_n263_3472.n6 a_n263_3472.t2 1.99806
R18782 a_n263_3472.n6 a_n263_3472.t1 1.99806
R18783 a_n263_3472.n4 a_n263_3472.t4 1.99806
R18784 a_n263_3472.n4 a_n263_3472.t3 1.99806
R18785 a_n263_3472.n5 a_n263_3472.t7 1.99806
R18786 a_n263_3472.n5 a_n263_3472.t5 1.99806
R18787 a_n263_3472.n2 a_n263_3472.t11 1.4923
R18788 a_n263_3472.n3 a_n263_3472.t8 1.4923
R18789 a_n263_3472.n8 a_n263_3472.t14 1.4923
R18790 a_n263_3472.n11 a_n263_3472.t12 1.4923
R18791 a_n263_3472.n0 a_n263_3472.n1 1.35826
R18792 a_21916_n6694.n20 a_21916_n6694.n19 25.8421
R18793 a_21916_n6694.n4 a_21916_n6694.n2 23.6976
R18794 a_21916_n6694.n5 a_21916_n6694.n1 22.4917
R18795 a_21916_n6694.n16 a_21916_n6694.t7 22.3385
R18796 a_21916_n6694.n12 a_21916_n6694.t16 18.9805
R18797 a_21916_n6694.n11 a_21916_n6694.t4 18.9805
R18798 a_21916_n6694.n7 a_21916_n6694.t15 18.9805
R18799 a_21916_n6694.n8 a_21916_n6694.t8 18.9805
R18800 a_21916_n6694.n1 a_21916_n6694.t21 18.6885
R18801 a_21916_n6694.n19 a_21916_n6694.t20 17.7395
R18802 a_21916_n6694.n4 a_21916_n6694.n3 17.1556
R18803 a_21916_n6694.n15 a_21916_n6694.t5 16.6445
R18804 a_21916_n6694.n12 a_21916_n6694.n11 16.5048
R18805 a_21916_n6694.n8 a_21916_n6694.n7 16.5048
R18806 a_21916_n6694.n15 a_21916_n6694.t14 15.4522
R18807 a_21916_n6694.n2 a_21916_n6694.t2 15.3305
R18808 a_21916_n6694.n18 a_21916_n6694.n14 15.3005
R18809 a_21916_n6694.n2 a_21916_n6694.t19 15.148
R18810 a_21916_n6694.n3 a_21916_n6694.t17 14.7222
R18811 a_21916_n6694.n3 a_21916_n6694.t18 14.6248
R18812 a_21916_n6694.n19 a_21916_n6694.t6 12.6782
R18813 a_21916_n6694.n1 a_21916_n6694.t9 11.8752
R18814 a_21916_n6694.n20 a_21916_n6694.n18 10.5305
R18815 a_21916_n6694.n21 a_21916_n6694.n20 10.4405
R18816 a_21916_n6694.n16 a_21916_n6694.t3 9.75817
R18817 a_21916_n6694.n17 a_21916_n6694.n15 9.01391
R18818 a_21916_n6694.n13 a_21916_n6694.t12 8.73617
R18819 a_21916_n6694.n10 a_21916_n6694.t10 8.73617
R18820 a_21916_n6694.n6 a_21916_n6694.t11 8.73617
R18821 a_21916_n6694.n9 a_21916_n6694.t13 8.73617
R18822 a_21916_n6694.n0 a_21916_n6694.n6 8.39376
R18823 a_21916_n6694.n0 a_21916_n6694.n10 8.3918
R18824 a_21916_n6694.n5 a_21916_n6694.n4 8.2805
R18825 a_21916_n6694.n17 a_21916_n6694.n16 8.01708
R18826 a_21916_n6694.n0 a_21916_n6694.n13 8.0005
R18827 a_21916_n6694.n0 a_21916_n6694.n9 8.0005
R18828 a_21916_n6694.n21 a_21916_n6694.t0 7.02774
R18829 a_21916_n6694.n13 a_21916_n6694.n12 6.0595
R18830 a_21916_n6694.n11 a_21916_n6694.n10 6.0595
R18831 a_21916_n6694.n7 a_21916_n6694.n6 6.0595
R18832 a_21916_n6694.n9 a_21916_n6694.n8 6.0595
R18833 a_21916_n6694.n14 a_21916_n6694.n0 5.41746
R18834 a_21916_n6694.n14 a_21916_n6694.n5 4.8605
R18835 a_21916_n6694.n18 a_21916_n6694.n17 4.8605
R18836 a_21916_n6694.t1 a_21916_n6694.n21 2.74964
R18837 a_23564_n452.t1 a_23564_n452.n3 50.3116
R18838 a_23564_n452.n2 a_23564_n452.t8 17.119
R18839 a_23564_n452.n0 a_23564_n452.t3 16.2065
R18840 a_23564_n452.n1 a_23564_n452.t5 16.2065
R18841 a_23564_n452.n3 a_23564_n452.t2 16.2065
R18842 a_23564_n452.n1 a_23564_n452.t7 13.1405
R18843 a_23564_n452.n3 a_23564_n452.t9 13.1405
R18844 a_23564_n452.n2 a_23564_n452.t6 12.228
R18845 a_23564_n452.n0 a_23564_n452.t4 12.228
R18846 a_23564_n452.n3 a_23564_n452.n1 10.5449
R18847 a_23564_n452.n3 a_23564_n452.n0 10.5449
R18848 a_23564_n452.t1 a_23564_n452.t0 9.70112
R18849 a_23564_n452.n0 a_23564_n452.n2 8.35614
R18850 a_24716_n5156.n0 a_24716_n5156.t5 29.2005
R18851 a_24716_n5156.n3 a_24716_n5156.n1 27.8386
R18852 a_24716_n5156.n3 a_24716_n5156.n2 24.9864
R18853 a_24716_n5156.n4 a_24716_n5156.n0 21.9516
R18854 a_24716_n5156.n2 a_24716_n5156.t2 20.1607
R18855 a_24716_n5156.n1 a_24716_n5156.t4 19.5523
R18856 a_24716_n5156.n0 a_24716_n5156.t7 12.1428
R18857 a_24716_n5156.n2 a_24716_n5156.t6 10.8288
R18858 a_24716_n5156.n1 a_24716_n5156.t3 9.79467
R18859 a_24716_n5156.n5 a_24716_n5156.n4 9.0005
R18860 a_24716_n5156.n5 a_24716_n5156.t0 8.32687
R18861 a_24716_n5156.n4 a_24716_n5156.n3 5.9405
R18862 a_24716_n5156.t1 a_24716_n5156.n5 4.54017
R18863 a_21804_n2273.n9 a_21804_n2273.n8 34.2905
R18864 a_21804_n2273.n0 a_21804_n2273.n5 19.9805
R18865 a_21804_n2273.n2 a_21804_n2273.t3 19.7105
R18866 a_21804_n2273.n3 a_21804_n2273.t2 19.7105
R18867 a_21804_n2273.n9 a_21804_n2273.n1 19.7105
R18868 a_21804_n2273.n5 a_21804_n2273.n4 17.9031
R18869 a_21804_n2273.t1 a_21804_n2273.n9 17.5055
R18870 a_21804_n2273.n7 a_21804_n2273.n0 17.2805
R18871 a_21804_n2273.n6 a_21804_n2273.t10 16.1822
R18872 a_21804_n2273.n8 a_21804_n2273.n2 15.8209
R18873 a_21804_n2273.n6 a_21804_n2273.t7 14.8925
R18874 a_21804_n2273.n2 a_21804_n2273.t12 13.3108
R18875 a_21804_n2273.n3 a_21804_n2273.t6 13.3108
R18876 a_21804_n2273.n7 a_21804_n2273.n6 12.6098
R18877 a_21804_n2273.n0 a_21804_n2273.t9 9.70587
R18878 a_21804_n2273.n5 a_21804_n2273.n3 8.7537
R18879 a_21804_n2273.n8 a_21804_n2273.n7 8.6405
R18880 a_21804_n2273.t1 a_21804_n2273.t0 8.3895
R18881 a_21804_n2273.n0 a_21804_n2273.t8 6.71423
R18882 a_21804_n2273.n1 a_21804_n2273.t13 6.71423
R18883 a_21804_n2273.n4 a_21804_n2273.t5 6.3005
R18884 a_21804_n2273.n4 a_21804_n2273.t4 5.6196
R18885 a_21804_n2273.n1 a_21804_n2273.t11 5.20587
R18886 a_22724_860.t7 a_22724_860.t5 161.001
R18887 a_22724_860.t4 a_22724_860.t6 104.147
R18888 a_22724_860.t5 a_22724_860.t2 33.5318
R18889 a_22724_860.t2 a_22724_860.t3 30.2103
R18890 a_22724_860.n0 a_22724_860.t7 17.9585
R18891 a_22724_860.t1 a_22724_860.t0 11.1158
R18892 a_22724_860.n0 a_22724_860.t4 8.07917
R18893 a_22724_860.t1 a_22724_860.n0 8.0005
R18894 a_23564_1116.t1 a_23564_1116.n3 53.3089
R18895 a_23564_1116.n2 a_23564_1116.t8 17.119
R18896 a_23564_1116.n0 a_23564_1116.t7 16.2065
R18897 a_23564_1116.n1 a_23564_1116.t9 16.2065
R18898 a_23564_1116.n3 a_23564_1116.t2 16.2065
R18899 a_23564_1116.n1 a_23564_1116.t5 13.1405
R18900 a_23564_1116.n3 a_23564_1116.t6 13.1405
R18901 a_23564_1116.n2 a_23564_1116.t4 12.228
R18902 a_23564_1116.n0 a_23564_1116.t3 12.228
R18903 a_23564_1116.n3 a_23564_1116.n1 10.5449
R18904 a_23564_1116.n3 a_23564_1116.n0 10.5449
R18905 a_23564_1116.t1 a_23564_1116.t0 8.3895
R18906 a_23564_1116.n0 a_23564_1116.n2 8.35614
R18907 a_23564_n14564.t1 a_23564_n14564.n3 36.9712
R18908 a_23564_n14564.n2 a_23564_n14564.t4 17.119
R18909 a_23564_n14564.n0 a_23564_n14564.t3 16.2065
R18910 a_23564_n14564.n1 a_23564_n14564.t5 16.2065
R18911 a_23564_n14564.n3 a_23564_n14564.t7 16.2065
R18912 a_23564_n14564.n1 a_23564_n14564.t9 13.1405
R18913 a_23564_n14564.n3 a_23564_n14564.t2 13.1405
R18914 a_23564_n14564.n2 a_23564_n14564.t8 12.228
R18915 a_23564_n14564.n0 a_23564_n14564.t6 12.228
R18916 a_23564_n14564.n3 a_23564_n14564.n1 10.5449
R18917 a_23564_n14564.n3 a_23564_n14564.n0 10.5449
R18918 a_23564_n14564.n0 a_23564_n14564.n2 8.35614
R18919 a_23564_n14564.t1 a_23564_n14564.t0 8.30886
R18920 a_28009_n1192.t1 a_28009_n1192.n0 54.9061
R18921 a_28009_n1192.n0 a_28009_n1192.t3 18.9805
R18922 a_28009_n1192.n0 a_28009_n1192.t2 11.4372
R18923 a_28009_n1192.t1 a_28009_n1192.t0 8.92356
R18924 a_21996_n12996.n10 a_21996_n12996.n9 40.4105
R18925 a_21996_n12996.n4 a_21996_n12996.n2 20.2983
R18926 a_21996_n12996.n1 a_21996_n12996.t10 17.484
R18927 a_21996_n12996.n7 a_21996_n12996.t11 17.484
R18928 a_21996_n12996.n5 a_21996_n12996.t5 17.484
R18929 a_21996_n12996.n3 a_21996_n12996.t6 17.484
R18930 a_21996_n12996.n2 a_21996_n12996.t12 17.484
R18931 a_21996_n12996.n4 a_21996_n12996.n3 17.4183
R18932 a_21996_n12996.n6 a_21996_n12996.n4 13.7705
R18933 a_21996_n12996.n9 a_21996_n12996.n1 12.7383
R18934 a_21996_n12996.n8 a_21996_n12996.n7 12.5636
R18935 a_21996_n12996.n6 a_21996_n12996.n5 12.5636
R18936 a_21996_n12996.n1 a_21996_n12996.t8 11.863
R18937 a_21996_n12996.n7 a_21996_n12996.t3 11.863
R18938 a_21996_n12996.n5 a_21996_n12996.t9 11.863
R18939 a_21996_n12996.n3 a_21996_n12996.t7 11.863
R18940 a_21996_n12996.n2 a_21996_n12996.t4 11.863
R18941 a_21996_n12996.n9 a_21996_n12996.n8 8.1455
R18942 a_21996_n12996.n10 a_21996_n12996.n0 6.83745
R18943 a_21996_n12996.n8 a_21996_n12996.n6 5.2205
R18944 a_21996_n12996.n0 a_21996_n12996.t1 3.37782
R18945 a_21996_n12996.n0 a_21996_n12996.t0 3.37782
R18946 a_21996_n12996.t2 a_21996_n12996.n10 3.03513
R18947 a_26060_n878.n0 a_26060_n878.n1 62.0943
R18948 a_26060_n878.n1 a_26060_n878.t2 18.141
R18949 a_26060_n878.n1 a_26060_n878.t3 11.863
R18950 a_26060_n878.n0 a_26060_n878.t1 8.56922
R18951 a_26060_n878.t0 a_26060_n878.n0 4.8813
R18952 a_25019_n3588.n5 a_25019_n3588.n3 29.1345
R18953 a_25019_n3588.n0 a_25019_n3588.t5 20.2215
R18954 a_25019_n3588.n2 a_25019_n3588.t9 20.2215
R18955 a_25019_n3588.n1 a_25019_n3588.n0 5.19536
R18956 a_25019_n3588.n3 a_25019_n3588.t6 18.6155
R18957 a_25019_n3588.n4 a_25019_n3588.t7 17.484
R18958 a_25019_n3588.n5 a_25019_n3588.n4 17.0878
R18959 a_25019_n3588.t1 a_25019_n3588.n6 16.2005
R18960 a_25019_n3588.n6 a_25019_n3588.n5 13.3205
R18961 a_25019_n3588.n3 a_25019_n3588.t4 11.8752
R18962 a_25019_n3588.n4 a_25019_n3588.t8 11.863
R18963 a_25019_n3588.n6 a_25019_n3588.n1 15.6414
R18964 a_25019_n3588.n1 a_25019_n3588.n2 5.09085
R18965 a_25019_n3588.n0 a_25019_n3588.t3 8.74833
R18966 a_25019_n3588.n2 a_25019_n3588.t2 8.74833
R18967 a_25019_n3588.t1 a_25019_n3588.t0 8.30886
R18968 XRST.n0 XRST.t2 19.7105
R18969 XRST.n0 XRST.t3 13.3108
R18970 XRST.n2 XRST.n0 8.9337
R18971 XRST.n1 XRST.t0 6.41334
R18972 XRST.n1 XRST.t1 5.50677
R18973 XRST.n2 XRST.n1 4.5005
R18974 XRST XRST.n2 3.84479
R18975 a_25836_n1236.n0 a_25836_n1236.n10 26.643
R18976 a_25836_n1236.n8 a_25836_n1236.t32 25.1125
R18977 a_25836_n1236.n7 a_25836_n1236.t23 25.1125
R18978 a_25836_n1236.n3 a_25836_n1236.n37 21.2539
R18979 a_25836_n1236.n35 a_25836_n1236.t20 20.1161
R18980 a_25836_n1236.n19 a_25836_n1236.n18 20.0683
R18981 a_25836_n1236.n19 a_25836_n1236.n17 19.2236
R18982 a_25836_n1236.n20 a_25836_n1236.t17 18.6885
R18983 a_25836_n1236.n35 a_25836_n1236.t41 18.2505
R18984 a_25836_n1236.n30 a_25836_n1236.t37 17.9585
R18985 a_25836_n1236.n27 a_25836_n1236.t36 17.9585
R18986 a_25836_n1236.n31 a_25836_n1236.t39 17.6787
R18987 a_25836_n1236.n26 a_25836_n1236.t8 17.6787
R18988 a_25836_n1236.n10 a_25836_n1236.t22 17.5205
R18989 a_25836_n1236.n17 a_25836_n1236.t10 17.484
R18990 a_25836_n1236.n12 a_25836_n1236.t38 17.4475
R18991 a_25836_n1236.n16 a_25836_n1236.t35 17.4475
R18992 a_25836_n1236.n13 a_25836_n1236.t12 17.4475
R18993 a_25836_n1236.n11 a_25836_n1236.t30 17.4475
R18994 a_25836_n1236.n34 a_25836_n1236.t25 17.3623
R18995 a_25836_n1236.n15 a_25836_n1236.n14 16.5048
R18996 a_25836_n1236.n31 a_25836_n1236.n30 16.5048
R18997 a_25836_n1236.n27 a_25836_n1236.n26 16.5048
R18998 a_25836_n1236.n12 a_25836_n1236.t26 16.3282
R18999 a_25836_n1236.n11 a_25836_n1236.t28 16.3282
R19000 a_25836_n1236.n18 a_25836_n1236.t29 15.4522
R19001 a_25836_n1236.n22 a_25836_n1236.t13 15.3305
R19002 a_25836_n1236.n18 a_25836_n1236.t9 15.1115
R19003 a_25836_n1236.n22 a_25836_n1236.t19 15.0872
R19004 a_25836_n1236.n15 a_25836_n1236.t18 14.7952
R19005 a_25836_n1236.n14 a_25836_n1236.t24 14.7952
R19006 a_25836_n1236.n34 a_25836_n1236.t16 14.6735
R19007 a_25836_n1236.n23 a_25836_n1236.n21 14.5805
R19008 a_25836_n1236.n23 a_25836_n1236.n22 12.8386
R19009 a_25836_n1236.n20 a_25836_n1236.t34 11.9603
R19010 a_25836_n1236.n17 a_25836_n1236.t14 11.863
R19011 a_25836_n1236.n10 a_25836_n1236.t40 11.5588
R19012 a_25836_n1236.n33 a_25836_n1236.n1 10.2605
R19013 a_25836_n1236.n9 a_25836_n1236.n7 9.94971
R19014 a_25836_n1236.n36 a_25836_n1236.n34 9.81008
R19015 a_25836_n1236.n2 a_25836_n1236.n12 9.01717
R19016 a_25836_n1236.n1 a_25836_n1236.n28 8.95618
R19017 a_25836_n1236.n21 a_25836_n1236.n20 8.90107
R19018 a_25836_n1236.n2 a_25836_n1236.n11 8.89383
R19019 a_25836_n1236.n29 a_25836_n1236.t27 8.80917
R19020 a_25836_n1236.n28 a_25836_n1236.t21 8.80917
R19021 a_25836_n1236.n8 a_25836_n1236.t15 8.73617
R19022 a_25836_n1236.n7 a_25836_n1236.t11 8.73617
R19023 a_25836_n1236.n37 a_25836_n1236.n33 8.4605
R19024 a_25836_n1236.n32 a_25836_n1236.t31 8.45633
R19025 a_25836_n1236.n25 a_25836_n1236.t33 8.45633
R19026 a_25836_n1236.n1 a_25836_n1236.n29 8.42898
R19027 a_25836_n1236.n1 a_25836_n1236.n25 8.4192
R19028 a_25836_n1236.n36 a_25836_n1236.n35 8.0005
R19029 a_25836_n1236.n9 a_25836_n1236.n8 8.0005
R19030 a_25836_n1236.n13 a_25836_n1236.n2 8.0005
R19031 a_25836_n1236.n2 a_25836_n1236.n16 8.0005
R19032 a_25836_n1236.n1 a_25836_n1236.n32 8.0005
R19033 a_25836_n1236.n3 a_25836_n1236.n5 7.10859
R19034 a_25836_n1236.n24 a_25836_n1236.n23 6.8405
R19035 a_25836_n1236.n3 a_25836_n1236.n6 6.32179
R19036 a_25836_n1236.n21 a_25836_n1236.n19 6.2555
R19037 a_25836_n1236.n0 a_25836_n1236.n2 6.04383
R19038 a_25836_n1236.n30 a_25836_n1236.n29 5.9865
R19039 a_25836_n1236.n28 a_25836_n1236.n27 5.9865
R19040 a_25836_n1236.n24 a_25836_n1236.n0 5.2205
R19041 a_25836_n1236.n0 a_25836_n1236.n9 5.1025
R19042 a_25836_n1236.n32 a_25836_n1236.n31 4.98883
R19043 a_25836_n1236.n26 a_25836_n1236.n25 4.98883
R19044 a_25836_n1236.n37 a_25836_n1236.n36 4.52892
R19045 a_25836_n1236.n3 a_25836_n1236.n4 3.40569
R19046 a_25836_n1236.n38 a_25836_n1236.n3 2.90888
R19047 a_25836_n1236.n33 a_25836_n1236.n24 2.7005
R19048 a_25836_n1236.n6 a_25836_n1236.t0 2.01032
R19049 a_25836_n1236.n6 a_25836_n1236.t2 2.01032
R19050 a_25836_n1236.n5 a_25836_n1236.t1 2.01032
R19051 a_25836_n1236.n5 a_25836_n1236.t3 2.01032
R19052 a_25836_n1236.n16 a_25836_n1236.n15 1.5335
R19053 a_25836_n1236.n14 a_25836_n1236.n13 1.5335
R19054 a_25836_n1236.n4 a_25836_n1236.t6 1.49844
R19055 a_25836_n1236.n4 a_25836_n1236.t4 1.49844
R19056 a_25836_n1236.t7 a_25836_n1236.n38 1.49844
R19057 a_25836_n1236.n38 a_25836_n1236.t5 1.49844
R19058 a_27337_1944.t1 a_27337_1944.n0 49.4957
R19059 a_27337_1944.n0 a_27337_1944.t2 17.5205
R19060 a_27337_1944.n0 a_27337_1944.t3 11.5588
R19061 a_27337_1944.t1 a_27337_1944.t0 8.92356
R19062 OUT[4] OUT[4].n14 19.5125
R19063 OUT[4].n3 OUT[4].n2 6.90733
R19064 OUT[4].n3 OUT[4].n1 6.3768
R19065 OUT[4].n12 OUT[4].n0 6.3768
R19066 OUT[4].n14 OUT[4].n13 6.3005
R19067 OUT[4].n9 OUT[4].n8 3.23472
R19068 OUT[4].n6 OUT[4].n5 3.21104
R19069 OUT[4].n9 OUT[4].n7 2.7042
R19070 OUT[4].n6 OUT[4].n4 2.7042
R19071 OUT[4].n7 OUT[4].t14 2.06607
R19072 OUT[4].n8 OUT[4].t13 2.06607
R19073 OUT[4].n5 OUT[4].t9 2.06607
R19074 OUT[4].n4 OUT[4].t11 2.06607
R19075 OUT[4].n13 OUT[4].t4 1.99806
R19076 OUT[4].n13 OUT[4].t1 1.99806
R19077 OUT[4].n2 OUT[4].t5 1.99806
R19078 OUT[4].n2 OUT[4].t2 1.99806
R19079 OUT[4].n1 OUT[4].t6 1.99806
R19080 OUT[4].n1 OUT[4].t0 1.99806
R19081 OUT[4].n0 OUT[4].t3 1.99806
R19082 OUT[4].n0 OUT[4].t7 1.99806
R19083 OUT[4].n7 OUT[4].t8 1.4923
R19084 OUT[4].n8 OUT[4].t10 1.4923
R19085 OUT[4].n5 OUT[4].t12 1.4923
R19086 OUT[4].n4 OUT[4].t15 1.4923
R19087 OUT[4].n14 OUT[4].n12 0.577837
R19088 OUT[4].n11 OUT[4].n3 0.189974
R19089 OUT[4].n10 OUT[4].n6 0.175763
R19090 OUT[4].n10 OUT[4].n9 0.166289
R19091 OUT[4].n12 OUT[4].n11 0.152079
R19092 OUT[4].n11 OUT[4].n10 0.145625
R19093 VIN VIN.t0 70.0209
R19094 a_22264_n1148.t1 a_22264_n1148.n0 66.3236
R19095 a_22264_n1148.n0 a_22264_n1148.t3 13.5573
R19096 a_22264_n1148.n0 a_22264_n1148.t2 11.0235
R19097 a_22264_n1148.t1 a_22264_n1148.t0 10.0058
R19098 a_34428_n452.n3 a_34428_n452.t3 29.2005
R19099 a_34428_n452.n4 a_34428_n452.n3 28.9716
R19100 a_34428_n452.n2 a_34428_n452.n0 23.6425
R19101 a_34428_n452.n1 a_34428_n452.t4 19.7105
R19102 a_34428_n452.n0 a_34428_n452.t5 17.2528
R19103 a_34428_n452.n2 a_34428_n452.n1 14.0209
R19104 a_34428_n452.n1 a_34428_n452.t7 13.3108
R19105 a_34428_n452.n0 a_34428_n452.t2 12.1672
R19106 a_34428_n452.n3 a_34428_n452.t6 12.1428
R19107 a_34428_n452.t1 a_34428_n452.t0 8.76859
R19108 a_34428_n452.n4 a_34428_n452.n2 7.5605
R19109 a_34428_n452.t1 a_34428_n452.n4 4.70222
R19110 a_23564_n3588.t1 a_23564_n3588.n3 46.6627
R19111 a_23564_n3588.n2 a_23564_n3588.t3 17.119
R19112 a_23564_n3588.n0 a_23564_n3588.t9 16.2065
R19113 a_23564_n3588.n1 a_23564_n3588.t8 16.2065
R19114 a_23564_n3588.n3 a_23564_n3588.t6 16.2065
R19115 a_23564_n3588.n1 a_23564_n3588.t7 13.1405
R19116 a_23564_n3588.n3 a_23564_n3588.t5 13.1405
R19117 a_23564_n3588.n2 a_23564_n3588.t2 12.228
R19118 a_23564_n3588.n0 a_23564_n3588.t4 12.228
R19119 a_23564_n3588.n3 a_23564_n3588.n1 10.5449
R19120 a_23564_n3588.n3 a_23564_n3588.n0 10.5449
R19121 a_23564_n3588.t1 a_23564_n3588.t0 9.70112
R19122 a_23564_n3588.n0 a_23564_n3588.n2 8.35614
R19123 a_29900_n10600.n3 a_29900_n10600.n4 32.8521
R19124 a_29900_n10600.n3 a_29900_n10600.n5 31.1127
R19125 a_29900_n10600.n0 a_29900_n10600.t9 20.2945
R19126 a_29900_n10600.n2 a_29900_n10600.t4 20.2945
R19127 a_29900_n10600.n1 a_29900_n10600.n0 5.17048
R19128 a_29900_n10600.n5 a_29900_n10600.t3 18.9805
R19129 a_29900_n10600.n4 a_29900_n10600.t5 18.6885
R19130 a_29900_n10600.n4 a_29900_n10600.t8 11.8752
R19131 a_29900_n10600.n5 a_29900_n10600.t2 11.4372
R19132 a_29900_n10600.n3 a_29900_n10600.n1 8.21661
R19133 a_29900_n10600.n1 a_29900_n10600.n2 5.11574
R19134 a_29900_n10600.n0 a_29900_n10600.t7 8.73617
R19135 a_29900_n10600.n2 a_29900_n10600.t6 8.73617
R19136 a_29900_n10600.t1 a_29900_n10600.t0 8.30886
R19137 a_29900_n10600.t1 a_29900_n10600.n3 7.1105
R19138 a_28852_n8292.n0 a_28852_n8292.n1 37.3822
R19139 a_28852_n8292.n1 a_28852_n8292.t3 17.4475
R19140 a_28852_n8292.n1 a_28852_n8292.t2 12.7755
R19141 a_28852_n8292.n0 a_28852_n8292.t1 8.31075
R19142 a_28852_n8292.t0 a_28852_n8292.n0 5.13976
R19143 a_25076_n4.n1 a_25076_n4.n0 58.1378
R19144 a_25076_n4.n0 a_25076_n4.t2 17.8003
R19145 a_25076_n4.n0 a_25076_n4.t3 14.7465
R19146 a_25076_n4.n1 a_25076_n4.t0 9.61569
R19147 a_25076_n4.t1 a_25076_n4.n1 4.52215
R19148 a_22892_n5156.n1 a_22892_n5156.n0 42.4705
R19149 a_22892_n5156.n0 a_22892_n5156.t4 17.484
R19150 a_22892_n5156.n0 a_22892_n5156.t3 11.863
R19151 a_22892_n5156.n1 a_22892_n5156.t1 6.58175
R19152 a_22892_n5156.t1 a_22892_n5156.t2 5.92991
R19153 a_22892_n5156.t0 a_22892_n5156.n1 5.70053
R19154 a_28940_n2406.n5 a_28940_n2406.n4 25.1646
R19155 a_28940_n2406.n3 a_28940_n2406.n2 20.9698
R19156 a_28940_n2406.n5 a_28940_n2406.n3 20.1605
R19157 a_28940_n2406.n0 a_28940_n2406.n5 19.4405
R19158 a_28940_n2406.n1 a_28940_n2406.t5 18.3235
R19159 a_28940_n2406.n2 a_28940_n2406.t7 18.3235
R19160 a_28940_n2406.n3 a_28940_n2406.n1 17.2494
R19161 a_28940_n2406.n4 a_28940_n2406.t2 17.119
R19162 a_28940_n2406.n1 a_28940_n2406.t4 12.7633
R19163 a_28940_n2406.n2 a_28940_n2406.t6 12.7633
R19164 a_28940_n2406.n4 a_28940_n2406.t3 12.7147
R19165 a_28940_n2406.n0 a_28940_n2406.t0 8.56922
R19166 a_28940_n2406.t1 a_28940_n2406.n0 4.8813
R19167 a_26172_n14564.t0 a_26172_n14564.n0 51.0033
R19168 a_26172_n14564.n0 a_26172_n14564.t2 18.141
R19169 a_26172_n14564.n0 a_26172_n14564.t3 11.863
R19170 a_26172_n14564.t0 a_26172_n14564.t1 9.23556
R19171 a_23703_n5156.n6 a_23703_n5156.n4 22.8155
R19172 a_23703_n5156.n1 a_23703_n5156.t7 18.3235
R19173 a_23703_n5156.n0 a_23703_n5156.t6 18.3235
R19174 a_23703_n5156.n5 a_23703_n5156.t8 18.2505
R19175 a_23703_n5156.n2 a_23703_n5156.t2 18.2505
R19176 a_23703_n5156.n3 a_23703_n5156.t9 18.2505
R19177 a_23703_n5156.n8 a_23703_n5156.n7 16.3805
R19178 a_23703_n5156.n4 a_23703_n5156.n3 14.7294
R19179 a_23703_n5156.n8 a_23703_n5156.n0 14.6816
R19180 a_23703_n5156.n7 a_23703_n5156.n1 12.9294
R19181 a_23703_n5156.n5 a_23703_n5156.t10 12.8242
R19182 a_23703_n5156.n2 a_23703_n5156.t3 12.8242
R19183 a_23703_n5156.n3 a_23703_n5156.t11 12.8242
R19184 a_23703_n5156.n1 a_23703_n5156.t4 12.7633
R19185 a_23703_n5156.n0 a_23703_n5156.t5 12.7633
R19186 a_23703_n5156.n6 a_23703_n5156.n5 12.7466
R19187 a_23703_n5156.n4 a_23703_n5156.n2 12.7466
R19188 a_23703_n5156.n9 a_23703_n5156.t0 6.92347
R19189 a_23703_n5156.n9 a_23703_n5156.n8 4.6355
R19190 a_23703_n5156.n7 a_23703_n5156.n6 3.9155
R19191 a_23703_n5156.t1 a_23703_n5156.n9 2.85249
R19192 a_29263_n3588.n0 a_29263_n3588.n1 40.1113
R19193 a_29263_n3588.n1 a_29263_n3588.t2 16.4012
R19194 a_29263_n3588.n1 a_29263_n3588.t3 14.6735
R19195 a_29263_n3588.n0 a_29263_n3588.t1 8.31075
R19196 a_29263_n3588.t0 a_29263_n3588.n0 5.13976
R19197 a_23999_n2320.n0 a_23999_n2320.n1 34.5269
R19198 a_23999_n2320.n2 a_23999_n2320.t5 29.2005
R19199 a_23999_n2320.n0 a_23999_n2320.n3 19.8281
R19200 a_23999_n2320.n1 a_23999_n2320.t6 19.7105
R19201 a_23999_n2320.n0 a_23999_n2320.n2 17.6316
R19202 a_23999_n2320.n3 a_23999_n2320.t4 16.3403
R19203 a_23999_n2320.n3 a_23999_n2320.t3 14.7465
R19204 a_23999_n2320.n1 a_23999_n2320.t2 13.3108
R19205 a_23999_n2320.n2 a_23999_n2320.t7 12.1428
R19206 a_23999_n2320.t1 a_23999_n2320.n0 11.7222
R19207 a_23999_n2320.t1 a_23999_n2320.t0 8.76859
R19208 a_25539_n407.n2 a_25539_n407.n0 37.8698
R19209 a_25539_n407.n1 a_25539_n407.t5 29.2005
R19210 a_25539_n407.n2 a_25539_n407.n1 21.0516
R19211 a_25539_n407.n0 a_25539_n407.t2 19.7105
R19212 a_25539_n407.n0 a_25539_n407.t4 13.3108
R19213 a_25539_n407.n1 a_25539_n407.t3 12.1428
R19214 a_25539_n407.t1 a_25539_n407.n2 10.2822
R19215 a_25539_n407.t1 a_25539_n407.t0 8.76859
R19216 a_27001_n4328.t1 a_27001_n4328.n0 46.7507
R19217 a_27001_n4328.n0 a_27001_n4328.t3 17.5205
R19218 a_27001_n4328.n0 a_27001_n4328.t2 11.5588
R19219 a_27001_n4328.t1 a_27001_n4328.t0 8.92356
R19220 a_24731_n3124.t0 a_24731_n3124.n2 38.0337
R19221 a_24731_n3124.n2 a_24731_n3124.n1 18.2371
R19222 a_24731_n3124.n0 a_24731_n3124.t3 17.7395
R19223 a_24731_n3124.n1 a_24731_n3124.t2 17.7395
R19224 a_24731_n3124.n2 a_24731_n3124.n0 17.3821
R19225 a_24731_n3124.n0 a_24731_n3124.t5 12.6782
R19226 a_24731_n3124.n1 a_24731_n3124.t4 12.6782
R19227 a_24731_n3124.t0 a_24731_n3124.t1 8.84645
R19228 a_33820_n452.t1 a_33820_n452.n0 34.5853
R19229 a_33820_n452.n0 a_33820_n452.t3 21.499
R19230 a_33820_n452.t1 a_33820_n452.t0 8.92356
R19231 a_33820_n452.n0 a_33820_n452.t2 8.69967
R19232 a_22276_n1572.t1 a_22276_n1572.n0 51.2292
R19233 a_22276_n1572.n0 a_22276_n1572.t2 19.7105
R19234 a_22276_n1572.n0 a_22276_n1572.t3 13.3108
R19235 a_22276_n1572.t1 a_22276_n1572.t0 9.70112
R19236 a_25795_n2716.t6 a_25795_n2716.t7 161.001
R19237 a_25795_n2716.t5 a_25795_n2716.t4 104.147
R19238 a_25795_n2716.t7 a_25795_n2716.t2 33.5318
R19239 a_25795_n2716.t2 a_25795_n2716.t3 30.2103
R19240 a_25795_n2716.n0 a_25795_n2716.t6 17.9585
R19241 a_25795_n2716.t1 a_25795_n2716.t0 11.1158
R19242 a_25795_n2716.n0 a_25795_n2716.t5 8.07917
R19243 a_25795_n2716.t1 a_25795_n2716.n0 8.0005
R19244 a_22668_n14864.n1 a_22668_n14864.n0 30.693
R19245 a_22668_n14864.n0 a_22668_n14864.t2 17.5205
R19246 a_22668_n14864.n0 a_22668_n14864.t3 11.5588
R19247 a_22668_n14864.n1 a_22668_n14864.t0 9.61569
R19248 a_22668_n14864.t1 a_22668_n14864.n1 4.52215
R19249 a_24716_1208.n2 a_24716_1208.n1 30.3851
R19250 a_24716_1208.n0 a_24716_1208.t5 29.2005
R19251 a_24716_1208.n1 a_24716_1208.t2 20.1607
R19252 a_24716_1208.n2 a_24716_1208.n0 19.2516
R19253 a_24716_1208.n0 a_24716_1208.t4 12.1428
R19254 a_24716_1208.n1 a_24716_1208.t3 10.8288
R19255 a_24716_1208.t1 a_24716_1208.n2 9.0005
R19256 a_24716_1208.t1 a_24716_1208.t0 8.44273
R19257 a_27225_n1572.t1 a_27225_n1572.n0 56.8183
R19258 a_27225_n1572.n0 a_27225_n1572.t2 18.9805
R19259 a_27225_n1572.n0 a_27225_n1572.t3 11.4372
R19260 a_27225_n1572.t1 a_27225_n1572.t0 8.92356
R19261 a_21692_n7508.n1 a_21692_n7508.n0 41.403
R19262 a_21692_n7508.n0 a_21692_n7508.t2 17.5205
R19263 a_21692_n7508.n0 a_21692_n7508.t3 11.5588
R19264 a_21692_n7508.n1 a_21692_n7508.t0 9.61569
R19265 a_21692_n7508.t1 a_21692_n7508.n1 4.52215
C0 a_41652_n3140 VDD 0.205948f
C1 a_22016_n10529 a_24233_n10252 0.020455f
C2 a_21604_n10116 a_23816_n10112 0.042802f
C3 a_21772_n9860 a_24684_n16432 0.033744f
C4 a_36192_1248 VDD 0.010384f
C5 a_32351_n7376 VDD 0.02509f
C6 a_21940_n11684 a_22352_n12097 0.536965f
C7 a_32424_n10512 VDD 0.363287f
C8 a_22772_n13648 VDD 0.299822f
C9 a_24315_n2759 a_23507_n2759 0.021748f
C10 a_46668_n14213 a_46580_n14116 0.285629f
C11 a_37844_n14116 a_38292_n14116 0.013276f
C12 a_39648_n2020 a_40196_n1884 0.239423f
C13 a_22500_n1976 a_23816_n704 0.022346f
C14 a_42188_n3237 a_42100_n3140 0.285629f
C15 a_46220_n3237 a_46668_n3237 0.012882f
C16 a_34872_1619 a_35849_n1192 0.014861f
C17 a_37844_n18820 VDD 0.215166f
C18 a_31324_n4372 a_24631_n3588 1.20173f
C19 a_27988_n17252 a_27988_n18440 0.05841f
C20 a_41204_n17252 a_41652_n17252 0.013276f
C21 a_46668_n4805 a_46580_n4708 0.285629f
C22 a_36588_n18917 a_36500_n18820 0.285629f
C23 a_31996_n20485 a_32444_n20485 0.013103f
C24 a_28435_n10599 a_30808_n10116 0.40326f
C25 a_29992_n11150 a_29744_n10980 0.370067f
C26 a_46468_n7464 VDD 0.209055f
C27 a_25573_n12167 a_25472_n14816 0.04547f
C28 a_44092_n10644 VDD 0.3211f
C29 a_23816_n13248 a_25237_n13735 0.015313f
C30 a_26563_n12212 a_27404_n14990 0.427305f
C31 a_22016_n13665 a_24128_n13248 0.277491f
C32 a_41764_n13736 VDD 0.206217f
C33 a_46556_n1669 a_46468_n1572 0.285629f
C34 a_27988_n4328 a_31412_n2276 0.044354f
C35 a_43556_n16872 VDD 0.209225f
C36 a_23844_n16872 a_23932_n16916 0.285629f
C37 a_22140_n16916 a_22588_n16916 0.012552f
C38 a_23484_n20052 VDD 0.318186f
C39 a_21604_n5412 a_22568_n5808 0.08126f
C40 a_22016_n5825 a_22364_n5808 0.401636f
C41 a_22052_n18440 a_21692_n18484 0.087174f
C42 a_35604_n17252 a_35716_n18440 0.026657f
C43 a_33812_n18820 a_34260_n18820 0.013276f
C44 a_47116_n18917 a_47476_n18820 0.087066f
C45 a_42157_n660 VDD 0.685388f
C46 a_40420_n9032 a_40060_n9076 0.087066f
C47 a_32444_n20485 a_32356_n20388 0.285629f
C48 a_25860_n9032 a_26266_n9240 0.026402f
C49 a_44004_n9032 a_44452_n9032 0.013276f
C50 a_25573_n12167 a_24965_n9860 0.048871f
C51 a_46468_n4328 VDD 0.209055f
C52 a_43725_908 VDD 0.702246f
C53 a_42636_n7941 VDD 0.313885f
C54 a_35804_n12212 a_36252_n12212 0.012552f
C55 a_25084_1564 OUT[1] 0.031891f
C56 a_35064_n11383 VDD 0.472952f
C57 a_27192_n14286 VDD 0.40616f
C58 a_33364_n15304 a_33812_n15304 0.013276f
C59 a_24403_n2414 a_23507_n2759 0.024286f
C60 a_43444_n14116 a_43556_n15304 0.026657f
C61 a_33452_n17349 VDD 0.320102f
C62 a_23564_n17700 a_24604_n17349 0.029576f
C63 a_32580_n16872 a_32220_n16916 0.087174f
C64 a_27572_860 a_28492_332 0.016589f
C65 a_37284_n20008 VDD 0.231657f
C66 a_42548_n17252 a_42660_n18440 0.026657f
C67 a_29892_n18440 a_30340_n18440 0.013276f
C68 a_46132_n4708 a_46020_n5896 0.026657f
C69 a_22444_n5156 a_22712_n7420 0.018497f
C70 a_42300_n7508 a_42748_n7508 0.012882f
C71 a_45572_n9032 a_45212_n9076 0.086905f
C72 a_43420_n20485 a_43780_n20388 0.087174f
C73 a_40060_n10644 a_40508_n10644 0.012882f
C74 a_44004_n10600 a_44092_n10644 0.285629f
C75 a_42660_n12168 a_42300_n12212 0.087066f
C76 a_41652_n10980 VDD 0.205948f
C77 a_37732_n13736 a_38180_n13736 0.013276f
C78 a_48012_n14213 VDD 0.343411f
C79 a_32020_n2276 a_31392_n2760 0.105654f
C80 a_24631_n3588 a_30408_n1104 0.036864f
C81 a_40652_n1572 a_45124_n1192 0.014911f
C82 a_37859_377 a_41684_n1976 0.116175f
C83 a_34260_n17252 VDD 0.205948f
C84 a_23564_n17700 a_28436_n17252 0.029641f
C85 a_39524_n16872 a_39972_n16872 0.013276f
C86 a_21604_n3844 a_22444_n5156 0.031349f
C87 a_43644_n705 a_45572_376 0.013789f
C88 a_45012_1564 a_45124_376 0.026657f
C89 a_47900_n20052 VDD 0.351088f
C90 a_40172_n5940 a_40620_n5940 0.013103f
C91 a_43668_n5896 a_43756_n5940 0.285629f
C92 a_42300_n7508 CLK 0.05218f
C93 a_23396_n20008 a_23484_n20052 0.285629f
C94 a_26980_n20008 a_27428_n20008 0.013276f
C95 a_40508_n7508 a_40396_n7941 0.026339f
C96 a_22712_n7420 a_26861_n8567 0.015774f
C97 a_44764_n1669 VDD 0.341707f
C98 a_23564_n8292 a_23564_n11428 1.65135f
C99 a_44340_n4708 VDD 0.214333f
C100 a_21772_n9860 a_24573_n12996 0.024554f
C101 a_37284_n9032 VDD 0.2329f
C102 a_47364_n12168 a_47452_n12212 0.285629f
C103 a_36700_n12212 a_36812_n12645 0.026339f
C104 a_45660_n12212 a_46108_n12212 0.012552f
C105 a_36612_n12168 VDD 0.215761f
C106 a_31664_n13292 a_31789_n14564 0.033441f
C107 a_37785_n364 a_38733_n727 0.016355f
C108 a_23708_n15216 VDD 0.012114f
C109 a_22164_n2760 a_27337_n3140 0.076442f
C110 a_40956_n15348 a_41404_n15348 0.012882f
C111 a_22820_n2804 a_25600_n5895 0.023713f
C112 a_23004_n2332 a_22588_n2020 0.059437f
C113 a_22140_n18484 VDD 0.296789f
C114 a_42300_n4372 a_42748_n4372 0.012552f
C115 a_23564_n17700 a_23396_n18440 0.035046f
C116 a_39056_820 a_39308_n452 0.031941f
C117 a_39056_820 a_38951_420 0.536965f
C118 a_38295_332 a_38847_464 0.119687f
C119 a_47228_n20485 VDD 0.329378f
C120 a_39972_n18440 a_40060_n18484 0.285629f
C121 a_23887_n5156 a_23564_n8292 0.033556f
C122 a_43556_n18440 a_44004_n18440 0.013276f
C123 a_38156_n7941 a_38604_n7941 0.013103f
C124 a_44340_n18820 a_44452_n20008 0.026657f
C125 a_23319_n2759 VDD 0.913643f
C126 a_40084_n5896 VDD 0.12475f
C127 a_25724_n14564 a_25559_n12548 0.010559f
C128 a_45212_n10644 a_45324_n11077 0.026339f
C129 a_29744_n10980 a_30296_n10980 0.361958f
C130 a_47452_n9076 VDD 0.313885f
C131 a_27744_n12908 a_28040_n12493 0.05539f
C132 a_41852_n12212 VDD 0.315469f
C133 a_29444_n708 a_29295_n1400 0.021163f
C134 a_41764_n15304 VDD 0.206217f
C135 a_45572_n2760 a_46020_n2760 0.013276f
C136 a_39164_n15348 a_39276_n15781 0.026339f
C137 a_32860_n2020 a_36520_n3868 0.024916f
C138 a_25759_1944 a_26383_1944 0.104193f
C139 a_36700_n18484 VDD 0.347096f
C140 a_28972_n17349 a_29420_n17349 0.013103f
C141 a_22444_n5156 a_24492_n5156 0.060108f
C142 a_22544_n4690 a_23479_n5156 0.03472f
C143 a_27988_n4328 a_26973_n8292 0.011848f
C144 a_47588_n20388 VDD 0.209676f
C145 a_45572_376 a_45660_332 0.285629f
C146 a_47900_n5940 a_48012_n6373 0.026339f
C147 a_45572_n18440 a_45212_n18484 0.086905f
C148 a_30215_n6265 a_30808_n6334 0.361958f
C149 a_33116_n20052 a_33564_n20052 0.012882f
C150 a_42636_n7941 a_42548_n7844 0.285629f
C151 a_37452_n3888 VDD 0.911043f
C152 a_25237_n10599 a_25412_n10600 0.26172f
C153 a_43532_n9509 a_43980_n9509 0.012882f
C154 a_23949_n6724 VDD 0.590784f
C155 a_36588_n9509 VDD 0.335291f
C156 a_37260_n12645 a_37708_n12645 0.012552f
C157 a_47476_n4 VDD 0.207033f
C158 a_22500_n15684 VDD 0.203482f
C159 a_37036_n15781 a_37484_n15781 0.012882f
C160 a_25237_n4327 a_25600_n5895 0.179957f
C161 a_47452_n18484 VDD 0.313885f
C162 a_28144_n4708 a_29612_n8292 1.05693f
C163 a_29420_n17349 a_29780_n17252 0.087174f
C164 a_27852_n18917 a_28300_n18917 0.012882f
C165 a_42188_n6373 a_42548_n6276 0.087066f
C166 a_24672_n11339 a_23816_n8544 0.02128f
C167 a_23479_n5156 a_21872_n9394 0.084499f
C168 a_22220_n9860 a_22016_n8961 0.023774f
C169 a_46132_n7844 a_46580_n7844 0.013276f
C170 a_40420_n20008 a_40060_n20052 0.087066f
C171 a_33588_n3461 VDD 1.75702f
C172 a_46668_n9509 a_47028_n9412 0.087066f
C173 a_47452_1900 VDD 0.336898f
C174 a_40308_n6276 VDD 0.211506f
C175 a_45324_n11077 a_45684_n10980 0.087066f
C176 a_37396_n10980 a_37844_n10980 0.013276f
C177 a_25573_n12167 a_25636_n14520 0.026027f
C178 a_25724_n14564 a_24233_n13388 0.032908f
C179 a_42996_n9412 VDD 0.205948f
C180 a_39500_n12645 a_39412_n12548 0.285629f
C181 a_34484_n12548 VDD 0.209253f
C182 a_46556_n1236 a_46556_n1669 0.05841f
C183 a_43980_n14213 a_44428_n14213 0.012882f
C184 a_35692_n14213 a_35604_n14116 0.285629f
C185 a_34708_n15684 VDD 0.205948f
C186 a_39276_n15781 a_39636_n15684 0.087066f
C187 a_22052_n15684 a_22052_n16872 0.05841f
C188 a_28153_1204 a_28048_1248 0.116059f
C189 a_42636_n18917 VDD 0.313885f
C190 a_23887_n5156 a_21604_n5412 0.013713f
C191 a_22544_n4690 a_22876_n5852 0.016366f
C192 a_29780_n17252 a_30228_n17252 0.013276f
C193 a_23479_n5156 a_22016_n5825 0.022168f
C194 a_40620_n17349 a_40532_n17252 0.285629f
C195 a_25612_n18917 a_25524_n18820 0.285629f
C196 a_47476_n6276 a_47924_n6276 0.013276f
C197 a_45572_n20008 a_45660_n20052 0.285629f
C198 a_46916_n20008 a_47364_n20008 0.013276f
C199 a_41204_n3140 VDD 0.227793f
C200 a_22364_n10512 a_22568_n10512 0.048436f
C201 a_21604_n10116 a_24233_n10252 0.019043f
C202 a_33048_n7420 VDD 0.361967f
C203 a_28300_n15348 a_33910_n12146 0.018161f
C204 a_32220_n10512 VDD 0.012291f
C205 a_41652_n12548 a_42100_n12548 0.013276f
C206 a_24128_n13248 VDD 0.024497f
C207 a_39648_n2020 a_37221_n3543 0.020182f
C208 a_46220_n14213 a_46580_n14116 0.087066f
C209 a_22500_n1976 a_24233_n844 0.017238f
C210 a_41740_n3237 a_42100_n3140 0.087066f
C211 a_41652_n15684 a_42100_n15684 0.013276f
C212 a_37396_n18820 VDD 0.212519f
C213 a_39972_n4708 a_40420_n4708 0.013276f
C214 a_46220_n4805 a_46580_n4708 0.087066f
C215 a_36140_n18917 a_36500_n18820 0.087066f
C216 a_22500_n18820 a_22948_n18820 0.013276f
C217 a_43444_n6276 a_43556_n7464 0.026657f
C218 a_46580_n7844 a_46468_n9032 0.026657f
C219 a_43444_n9412 a_43556_n10600 0.026657f
C220 a_46020_n7464 VDD 0.210736f
C221 a_42100_n10980 a_42212_n12168 0.026657f
C222 a_27281_n16854 a_27700_n14116 0.026091f
C223 a_43644_n10644 VDD 0.319164f
C224 a_24684_n16432 a_23564_n20836 0.010901f
C225 a_24233_n13388 a_25237_n13735 0.116758f
C226 a_41316_n13736 VDD 0.206217f
C227 a_32860_n2020 a_32020_n2276 0.049736f
C228 a_35604_n14116 a_35604_n15304 0.05841f
C229 a_27988_n4328 a_30555_n2729 0.463854f
C230 a_46108_n1669 a_46468_n1572 0.087174f
C231 a_43108_n16872 VDD 0.206217f
C232 a_37859_377 a_39556_n4 0.602643f
C233 a_23844_n16872 a_23484_n16916 0.086742f
C234 a_23036_n20052 VDD 0.315749f
C235 a_43833_1204 a_43644_n705 0.119778f
C236 a_22016_n5825 a_22876_n5852 0.882105f
C237 a_38180_n4708 a_38403_n5503 0.018983f
C238 a_21604_n5412 a_22364_n5808 0.011851f
C239 a_21604_n18440 a_21692_n18484 0.285629f
C240 a_24740_n18440 a_25188_n18440 0.013276f
C241 a_39076_n7464 a_39524_n7464 0.013276f
C242 a_22052_n6980 a_23564_n8292 0.128259f
C243 a_47116_n18917 a_47028_n18820 0.285629f
C244 a_41533_n727 VDD 0.586417f
C245 a_42972_n20485 a_43420_n20485 0.013103f
C246 a_39972_n9032 a_40060_n9076 0.285629f
C247 a_25860_n9032 a_25642_n9816 0.05829f
C248 a_31996_n20485 a_32356_n20388 0.087174f
C249 a_21872_n9394 a_21892_n9816 0.58475f
C250 a_46020_n4328 VDD 0.210736f
C251 a_43101_841 VDD 0.587175f
C252 a_42188_n7941 VDD 0.313885f
C253 a_30555_n13780 a_31455_n13648 0.116059f
C254 a_26944_n14116 VDD 0.804302f
C255 a_32556_n17349 VDD 0.338774f
C256 a_35268_n16872 a_35716_n16872 0.013276f
C257 a_32132_n16872 a_32220_n16916 0.285629f
C258 a_43892_n3140 a_44004_n4328 0.026657f
C259 a_36700_n20052 VDD 0.359864f
C260 a_22444_n5156 a_22464_n7393 0.015791f
C261 a_44340_n18820 a_44788_n18820 0.013276f
C262 a_25972_n6276 a_25573_n12167 0.072269f
C263 a_43420_n20485 a_43332_n20388 0.285629f
C264 a_25831_n11428 a_22220_n12996 0.037719f
C265 a_45124_n9032 a_45212_n9076 0.285629f
C266 a_46468_n9032 a_46916_n9032 0.013276f
C267 a_28548_n5112 VDD 0.020878f
C268 a_44004_n10600 a_43644_n10644 0.087066f
C269 a_42212_n12168 a_42300_n12212 0.285629f
C270 a_37820_n12212 a_38268_n12212 0.012882f
C271 a_41204_n10980 VDD 0.226701f
C272 a_44540_332 a_44509_n452 0.041366f
C273 a_47564_n14213 VDD 0.315469f
C274 a_32020_n2276 a_31412_n2276 0.10673f
C275 a_37732_n15304 a_38180_n15304 0.013276f
C276 a_33812_n17252 VDD 0.205948f
C277 a_39524_n4328 a_39972_n4328 0.013276f
C278 a_23564_n17700 a_27988_n17252 0.017768f
C279 a_21604_n3844 a_21604_n5067 0.029777f
C280 a_43644_n705 a_45124_376 0.033864f
C281 a_47452_n20052 VDD 0.328902f
C282 a_36612_n18440 a_36700_n18484 0.285629f
C283 a_32668_n18484 a_33116_n18484 0.012882f
C284 a_43668_n5896 a_43308_n5940 0.086742f
C285 a_41852_n7508 CLK 0.020312f
C286 a_22712_n7420 a_26531_n8639 0.213814f
C287 a_23396_n20008 a_23036_n20052 0.087066f
C288 a_44316_n1669 VDD 0.302649f
C289 a_43332_n20388 a_43780_n20388 0.013276f
C290 a_39612_n9076 a_39724_n9509 0.026339f
C291 a_43892_n4708 VDD 0.212278f
C292 a_47452_n10644 a_47900_n10644 0.012001f
C293 a_21772_n9860 a_23949_n12996 0.012408f
C294 a_47364_n12168 a_47004_n12212 0.086742f
C295 a_36164_n12168 VDD 0.208761f
C296 a_40508_n13780 a_40956_n13780 0.012882f
C297 a_44452_n13736 a_44540_n13780 0.285629f
C298 a_31664_n13292 a_28752_n15348 0.030229f
C299 a_21604_n708 a_22588_n2020 0.031746f
C300 a_24220_n15260 VDD 0.259213f
C301 a_41540_n2760 a_41988_n2760 0.013276f
C302 a_27988_n20388 a_28568_n16066 0.024784f
C303 a_28736_1944 a_28454_n2424 0.049874f
C304 a_21692_n18484 VDD 0.300735f
C305 a_34460_n16916 a_34348_n17349 0.026339f
C306 a_42300_n16916 a_42748_n16916 0.012882f
C307 a_37947_332 a_38847_464 0.116059f
C308 a_46780_n20485 VDD 0.33079f
C309 a_39972_n18440 a_39612_n18484 0.087066f
C310 a_29892_n20008 a_30340_n20008 0.013276f
C311 a_22672_n2759 VDD 0.595614f
C312 a_28435_n10599 a_32854_n12168 0.025446f
C313 a_29744_n10980 a_30092_n10980 0.401636f
C314 OUT[0] OUT[1] 0.026583f
C315 VDD OUT[4] 0.926684f
C316 a_47004_n9076 VDD 0.313885f
C317 a_43196_n12212 a_43084_n12645 0.026339f
C318 a_26983_n12728 a_28040_n12493 0.056721f
C319 a_25559_n12548 a_25132_n16432 0.239487f
C320 a_27281_n16854 a_27709_n16132 0.036873f
C321 a_41404_n12212 VDD 0.315469f
C322 a_41316_n15304 VDD 0.206217f
C323 a_21692_n15781 a_22140_n15781 0.012552f
C324 a_22052_1944 a_26607_1966 0.033638f
C325 a_36252_n18484 VDD 0.315469f
C326 a_41404_n16916 a_41292_n17349 0.026339f
C327 a_22444_n5156 a_23887_n5156 0.034896f
C328 a_22544_n4690 a_22788_n4708 0.015023f
C329 a_34068_n4 a_34272_n4 0.033243f
C330 a_46573_841 a_47197_908 0.104193f
C331 a_45572_376 a_45212_332 0.086742f
C332 a_47140_n20388 VDD 0.203482f
C333 a_30320_n6636 a_30616_n6221 0.05539f
C334 a_45124_n18440 a_45212_n18484 0.285629f
C335 a_46468_n18440 a_46916_n18440 0.013276f
C336 a_35804_n18484 a_35692_n18917 0.026339f
C337 a_23564_n8292 a_24128_n8544 0.049334f
C338 a_26973_n8292 a_26861_n8567 0.026651f
C339 a_42188_n7941 a_42548_n7844 0.087066f
C340 a_33188_n2672 VDD 0.299361f
C341 a_25237_n10599 a_23816_n10112 0.014425f
C342 a_23564_n8292 a_22352_n12097 0.023193f
C343 a_42188_n11077 a_42636_n11077 0.012882f
C344 a_34392_n9815 VDD 0.529151f
C345 a_46108_n13780 a_46220_n14213 0.026339f
C346 a_24578_n2020 a_25647_n1976 0.014406f
C347 a_22052_n15684 VDD 0.203482f
C348 a_27988_n4328 a_23479_n5156 0.051533f
C349 a_27672_n3543 a_27932_n3543 0.508765f
C350 a_22052_1944 a_29332_1243 0.067456f
C351 a_39748_2475 a_40196_1944 0.197353f
C352 a_47004_n18484 VDD 0.313885f
C353 a_45660_n4372 a_45772_n4805 0.026339f
C354 a_39724_n17349 a_40172_n17349 0.012882f
C355 a_29420_n17349 a_29332_n17252 0.285629f
C356 a_27988_n4328 a_29532_n10311 0.06619f
C357 a_22220_n9860 a_21604_n8548 0.037782f
C358 a_24672_n11339 a_24233_n8684 0.049566f
C359 a_42748_n18484 a_42636_n18917 0.026339f
C360 a_42188_n6373 a_42100_n6276 0.285629f
C361 a_47116_n6373 a_47564_n6373 0.012882f
C362 a_23479_n5156 a_27485_n8500 0.03405f
C363 a_39972_n20008 a_40060_n20052 0.285629f
C364 a_43556_n20008 a_44004_n20008 0.013276f
C365 a_46668_n9509 a_46580_n9412 0.285629f
C366 a_38740_n9412 a_39188_n9412 0.013276f
C367 a_29992_n11150 a_28435_n10599 0.578321f
C368 a_47364_1944 VDD 0.169751f
C369 a_39860_n6276 VDD 0.208018f
C370 a_45324_n11077 a_45236_n10980 0.285629f
C371 a_42548_n9412 VDD 0.205948f
C372 a_26983_n12728 a_26470_n13736 0.031936f
C373 a_39052_n12645 a_39412_n12548 0.086742f
C374 a_34036_n12548 VDD 0.123349f
C375 a_42524_n20485 CLK 0.022624f
C376 a_35244_n14213 a_35604_n14116 0.087066f
C377 a_34260_n15684 VDD 0.205948f
C378 a_47564_n15781 a_48012_n15781 0.012882f
C379 a_39276_n15781 a_39188_n15684 0.285629f
C380 a_27736_1248 a_28048_1248 0.119687f
C381 a_42188_n18917 VDD 0.313885f
C382 a_41292_n4805 a_41740_n4805 0.012882f
C383 a_40172_n17349 a_40532_n17252 0.086635f
C384 a_22544_n4690 a_22264_n5852 0.05466f
C385 a_38380_n18917 a_38828_n18917 0.012882f
C386 a_24828_n18917 a_25524_n18820 0.012267f
C387 a_45572_n20008 a_45212_n20052 0.086905f
C388 a_39412_n7844 a_39524_n9032 0.026657f
C389 a_40308_n3140 VDD 0.212206f
C390 a_22876_n10556 a_22568_n10512 0.934191f
C391 a_24965_n9860 a_24964_n14116 0.041494f
C392 a_41204_1243 VDD 1.80642f
C393 a_32455_n7420 VDD 0.803631f
C394 a_32732_n10556 VDD 0.248025f
C395 a_22500_n1976 a_28352_n320 0.020124f
C396 a_24315_n2759 a_24403_n2414 0.198709f
C397 a_21916_n1975 a_22672_n2759 0.01027f
C398 a_37396_n14116 a_37844_n14116 0.013276f
C399 a_46220_n14213 a_46132_n14116 0.285629f
C400 a_32636_n2020 a_34248_n3310 0.010205f
C401 a_27932_n3543 a_28144_n4708 0.604184f
C402 a_41740_n3237 a_41652_n3140 0.285629f
C403 a_45772_n3237 a_46220_n3237 0.012882f
C404 a_31324_n4372 a_31787_n3969 0.026638f
C405 a_28736_1944 a_24631_n3588 0.034092f
C406 a_35064_1506 a_35849_n1192 0.054548f
C407 a_34872_1619 a_35324_1564 0.026665f
C408 a_36948_n18820 VDD 0.213047f
C409 a_46220_n4805 a_46132_n4708 0.285629f
C410 a_24672_n11339 a_24965_n9860 0.066228f
C411 a_23479_n5156 a_26470_n9322 0.031926f
C412 a_36140_n18917 a_36052_n18820 0.285629f
C413 a_22016_n1121 VDD 0.796483f
C414 a_31548_n20485 a_31996_n20485 0.013103f
C415 a_28435_n10599 a_28247_n10599 0.26222f
C416 a_23004_n2332 VDD 0.791093f
C417 a_45572_n7464 VDD 0.213324f
C418 a_28121_n10980 a_27639_n12537 0.090956f
C419 a_27281_n16854 a_27496_n14116 0.033165f
C420 a_43196_n10644 VDD 0.316157f
C421 a_24233_n13388 a_23816_n13248 0.633318f
C422 a_40868_n13736 VDD 0.208618f
C423 a_46108_n1669 a_46020_n1572 0.285629f
C424 a_32636_n2020 a_32020_n2276 0.035638f
C425 a_42660_n16872 VDD 0.206217f
C426 a_23396_n16872 a_23484_n16916 0.285629f
C427 a_21692_n16916 a_22140_n16916 0.012552f
C428 a_37859_377 a_38996_n408 0.02038f
C429 a_37859_377 a_39544_420 0.037993f
C430 a_43416_1248 a_43644_n705 0.018961f
C431 a_22588_n20052 VDD 0.312663f
C432 a_22220_n9860 a_24573_n6724 0.06233f
C433 a_22016_n5825 a_22264_n5852 0.370731f
C434 a_21604_n5412 a_22876_n5852 0.05539f
C435 a_35156_n17252 a_35268_n18440 0.026657f
C436 a_46668_n18917 a_47028_n18820 0.087066f
C437 a_33364_n18820 a_33812_n18820 0.013276f
C438 a_29123_n6679 a_29532_n10311 0.031633f
C439 a_41203_n799 VDD 0.323102f
C440 a_31996_n20485 a_31908_n20388 0.285629f
C441 a_25860_n9032 a_25237_n10599 0.033313f
C442 a_43556_n9032 a_44004_n9032 0.013276f
C443 a_39972_n9032 a_39612_n9076 0.087066f
C444 a_45572_n4328 VDD 0.213324f
C445 a_25020_n11383 a_31856_n11296 0.012341f
C446 a_22264_n8988 a_22264_n13692 0.03134f
C447 a_42771_769 VDD 0.321307f
C448 a_21604_n10116 a_23564_n11428 0.067103f
C449 a_41740_n7941 VDD 0.313885f
C450 a_35356_n12212 a_35804_n12212 0.012552f
C451 a_31324_n4372 OUT[1] 0.034708f
C452 a_42996_n14116 a_43108_n15304 0.026657f
C453 a_32916_n15304 a_33364_n15304 0.013276f
C454 a_32108_n17349 VDD 0.320587f
C455 a_32132_n16872 a_31772_n16916 0.087174f
C456 a_36252_n20052 VDD 0.296789f
C457 a_22444_n5156 a_22052_n6980 0.01122f
C458 a_45684_n4708 a_45572_n5896 0.026657f
C459 a_36773_n5468 a_38733_n5431 0.016464f
C460 a_45772_n101 a_45684_n4 0.285629f
C461 a_29444_n18440 a_29892_n18440 0.013276f
C462 a_42100_n17252 a_42212_n18440 0.026657f
C463 a_41852_n7508 a_42300_n7508 0.012882f
C464 a_31908_n20388 a_32356_n20388 0.013276f
C465 a_42972_n20485 a_43332_n20388 0.087174f
C466 a_43556_n10600 a_43644_n10644 0.285629f
C467 a_39612_n10644 a_40060_n10644 0.012882f
C468 a_28009_n12168 a_28232_n12606 0.013122f
C469 a_42212_n12168 a_41852_n12212 0.087066f
C470 a_40532_n10980 VDD 0.213111f
C471 a_37284_n13736 a_37732_n13736 0.013276f
C472 a_31076_376 a_34068_n4 0.044334f
C473 a_47116_n14213 VDD 0.315469f
C474 a_31292_n2804 a_31412_n2276 0.406528f
C475 a_24631_n3588 a_30716_n1148 0.036743f
C476 a_33364_n17252 VDD 0.227793f
C477 a_23564_n17700 a_24516_n17252 0.055338f
C478 a_39076_n16872 a_39524_n16872 0.013276f
C479 a_47004_n20052 VDD 0.328902f
C480 a_43644_n705 a_44540_332 0.044936f
C481 a_43220_n5896 a_43308_n5940 0.285629f
C482 a_36612_n18440 a_36252_n18484 0.086635f
C483 a_41404_n7508 CLK 0.010246f
C484 a_26532_n20008 a_26980_n20008 0.013276f
C485 a_22712_n7420 a_23816_n8544 0.02693f
C486 a_40060_n7508 a_39948_n7941 0.026339f
C487 a_22948_n20008 a_23036_n20052 0.285629f
C488 a_43868_n1669 VDD 0.316035f
C489 a_43444_n4708 VDD 0.210872f
C490 a_21772_n9860 a_22264_n13692 0.034742f
C491 a_36252_n12212 a_36364_n12645 0.026339f
C492 a_46916_n12168 a_47004_n12212 0.285629f
C493 a_45212_n12212 a_45660_n12212 0.012552f
C494 a_35716_n12168 VDD 0.209244f
C495 a_21604_n708 a_21828_n1931 0.030334f
C496 a_44452_n13736 a_44092_n13780 0.086635f
C497 a_23608_n15260 VDD 0.578921f
C498 a_40508_n15348 a_40956_n15348 0.012882f
C499 a_27988_n20388 a_27709_n16132 0.028739f
C500 a_44452_n15304 a_44540_n15348 0.285629f
C501 a_22820_n2804 a_27337_n3140 0.012086f
C502 a_28736_1944 a_27452_n2716 0.823229f
C503 a_23004_n2332 a_21916_n1975 0.037863f
C504 a_28436_n18440 VDD 0.208933f
C505 a_28144_n4708 a_27414_n5112 0.239647f
C506 a_41852_n4372 a_42300_n4372 0.013103f
C507 a_38295_332 a_38951_420 0.510371f
C508 a_46332_n20485 VDD 0.333257f
C509 a_39524_n18440 a_39612_n18484 0.285629f
C510 a_43108_n18440 a_43556_n18440 0.013276f
C511 a_43892_n18820 a_44004_n20008 0.026657f
C512 a_37708_n7941 a_38156_n7941 0.013103f
C513 a_25139_n2704 VDD 0.256232f
C514 a_35568_n4 a_36120_n4 0.361958f
C515 a_39357_n5364 VDD 0.701947f
C516 a_29332_n11301 a_31961_n11340 0.019043f
C517 a_29744_n10980 a_30604_n11029 0.882105f
C518 a_46556_n9076 VDD 0.31705f
C519 a_27281_n16854 a_27085_n16132 0.055596f
C520 a_26983_n12728 a_27535_n12493 0.119687f
C521 a_24964_n14116 a_25636_n14520 0.010692f
C522 a_27744_n12908 a_28232_n12606 0.08126f
C523 a_40956_n12212 VDD 0.330158f
C524 a_26239_n12996 a_26755_n16132 0.214233f
C525 a_40868_n15304 VDD 0.208618f
C526 a_45124_n2760 a_45572_n2760 0.013276f
C527 a_38716_n15348 a_38828_n15781 0.026339f
C528 a_22052_1944 a_26383_1944 0.029599f
C529 a_35804_n18484 VDD 0.315469f
C530 a_22444_n5156 a_23479_n5156 0.084748f
C531 a_28524_n17349 a_28972_n17349 0.013103f
C532 a_46692_n20388 VDD 0.205569f
C533 a_45124_376 a_45212_332 0.285629f
C534 a_47452_n5940 a_47564_n6373 0.026339f
C535 a_29559_n6456 a_30616_n6221 0.056721f
C536 a_29612_n8292 a_29476_n6980 0.070835f
C537 a_32668_n20052 a_33116_n20052 0.012882f
C538 a_36612_n20008 a_36700_n20052 0.285629f
C539 a_42188_n7941 a_42100_n7844 0.285629f
C540 a_22712_n7420 a_25237_n10599 0.058291f
C541 a_23564_n8292 a_21940_n11684 0.01222f
C542 a_43084_n9509 a_43532_n9509 0.012882f
C543 a_24965_n9860 a_23816_n10112 0.048625f
C544 a_25237_n10599 a_24233_n10252 0.109494f
C545 a_32581_n9860 a_25020_n11383 0.510166f
C546 a_21812_n6643 VDD 0.837465f
C547 a_33494_n9860 VDD 0.596434f
C548 a_36812_n12645 a_37260_n12645 0.013103f
C549 a_24578_n2020 a_24315_n2759 0.488337f
C550 a_21604_n15684 VDD 0.221763f
C551 a_36588_n15781 a_37036_n15781 0.012882f
C552 a_47900_n15348 a_48012_n15781 0.026339f
C553 a_46556_n18484 VDD 0.31705f
C554 a_37859_377 a_40196_1944 0.042682f
C555 a_28972_n17349 a_29332_n17252 0.087174f
C556 a_27190_n5112 a_27414_n5112 0.75472f
C557 a_23479_n5156 a_26861_n8567 0.069067f
C558 a_27404_n18917 a_27852_n18917 0.012882f
C559 a_41740_n6373 a_42100_n6276 0.087066f
C560 a_39972_n20008 a_39612_n20052 0.087066f
C561 a_45684_n7844 a_46132_n7844 0.013276f
C562 a_25600_n5895 VDD 0.337005f
C563 a_46220_n9509 a_46580_n9412 0.087066f
C564 a_28437_n13705 a_28492_n12548 0.017864f
C565 a_36948_n10980 a_37396_n10980 0.013276f
C566 a_44876_n11077 a_45236_n10980 0.087066f
C567 a_42100_n9412 VDD 0.205948f
C568 a_39052_n12645 a_38964_n12548 0.285629f
C569 a_26563_n12212 a_27496_n14116 0.049352f
C570 a_25831_n12996 a_27526_n13714 0.295971f
C571 a_42076_n20485 CLK 0.029774f
C572 a_35244_n14213 a_35156_n14116 0.285629f
C573 a_43532_n14213 a_43980_n14213 0.012882f
C574 a_46108_n1236 a_46108_n1669 0.05841f
C575 a_33812_n15684 VDD 0.205948f
C576 a_21604_n15684 a_21604_n16872 0.05841f
C577 a_38828_n15781 a_39188_n15684 0.087066f
C578 a_36217_n3500 a_36112_n3456 0.116059f
C579 a_41740_n18917 VDD 0.313885f
C580 a_27736_1248 a_28153_1204 0.633318f
C581 a_29332_n17252 a_29780_n17252 0.013276f
C582 a_40172_n17349 a_40084_n17252 0.285629f
C583 a_22544_n4690 a_22016_n5825 0.040712f
C584 a_24828_n18917 a_24740_n18820 0.285629f
C585 a_47028_n6276 a_47476_n6276 0.013276f
C586 a_45124_n20008 a_45212_n20052 0.285629f
C587 a_46468_n20008 a_46916_n20008 0.013276f
C588 a_39860_n3140 VDD 0.208996f
C589 a_22016_n10529 a_22568_n10512 0.361958f
C590 a_32560_n7020 VDD 1.82053f
C591 a_31872_n10529 VDD 0.808271f
C592 a_41204_n12548 a_41652_n12548 0.013276f
C593 a_28736_1944 a_28456_n364 0.099936f
C594 a_42436_n20388 CLK 0.049487f
C595 a_27526_n13714 VDD 0.305943f
C596 a_45772_n14213 a_46132_n14116 0.087066f
C597 a_32636_n2020 a_34953_n1572 0.293584f
C598 a_41292_n3237 a_41652_n3140 0.087066f
C599 a_25600_n5895 a_26271_n4306 0.012786f
C600 a_41204_n15684 a_41652_n15684 0.013276f
C601 a_24628_1252 a_23136_447 0.035264f
C602 a_34471_1575 a_35849_n1192 0.400514f
C603 a_36500_n18820 VDD 0.208341f
C604 a_45772_n4805 a_46132_n4708 0.087066f
C605 a_39524_n4708 a_39972_n4708 0.013276f
C606 a_22052_n18820 a_22500_n18820 0.013276f
C607 a_35692_n18917 a_36052_n18820 0.087066f
C608 a_42996_n6276 a_43108_n7464 0.026657f
C609 a_24672_n11339 a_24573_n9860 0.066279f
C610 a_23479_n5156 a_26266_n9240 0.010349f
C611 a_21604_n708 VDD 1.82611f
C612 a_46132_n7844 a_46020_n9032 0.026657f
C613 a_28435_n10599 a_31460_n10116 0.044783f
C614 a_42996_n9412 a_43108_n10600 0.026657f
C615 a_45124_n7464 VDD 0.26277f
C616 a_41652_n10980 a_41764_n12168 0.026657f
C617 a_42748_n10644 VDD 0.315469f
C618 a_40420_n13736 VDD 0.206217f
C619 a_45660_n1669 a_46020_n1572 0.087174f
C620 a_35156_n14116 a_35156_n15304 0.05841f
C621 a_42212_n16872 VDD 0.206217f
C622 a_37859_377 a_39308_n452 0.286354f
C623 a_23396_n16872 a_23036_n16916 0.086742f
C624 a_47476_n3140 a_47924_n3140 0.013276f
C625 a_45100_1467 a_40652_n1572 0.048612f
C626 a_22140_n20052 VDD 0.312663f
C627 a_37859_377 a_38951_420 0.041271f
C628 a_24292_n18440 a_24740_n18440 0.013276f
C629 a_21604_n5412 a_22264_n5852 0.102497f
C630 a_38628_n7464 a_39076_n7464 0.013276f
C631 a_46668_n18917 a_46580_n18820 0.285629f
C632 a_39357_n660 VDD 0.731372f
C633 a_25412_n8501 a_25237_n10599 0.028848f
C634 a_31548_n20485 a_31908_n20388 0.087174f
C635 a_42524_n20485 a_42972_n20485 0.013103f
C636 a_39524_n9032 a_39612_n9076 0.285629f
C637 a_45124_n4328 VDD 0.26277f
C638 a_25020_n11383 a_31961_n11340 0.03245f
C639 a_32581_n9860 a_33572_n10980 0.015229f
C640 a_40776_770 VDD 0.40948f
C641 a_46580_n4 a_47028_n4 0.013276f
C642 a_41292_n7941 VDD 0.320102f
C643 a_31856_n11296 VDD 0.026192f
C644 a_30555_n13780 a_31559_n13692 0.020455f
C645 a_22164_n2760 a_23507_n2759 0.172055f
C646 a_28736_1944 a_28671_n1976 0.050987f
C647 a_35849_n1192 a_35119_n1170 0.234051f
C648 a_31660_n17349 VDD 0.329535f
C649 a_25237_n4327 a_32132_n4708 0.135609f
C650 a_43444_n3140 a_43556_n4328 0.026657f
C651 a_31684_n16872 a_31772_n16916 0.285629f
C652 a_34820_n16872 a_35268_n16872 0.013276f
C653 a_35804_n20052 VDD 0.296789f
C654 a_45324_n101 a_45684_n4 0.086905f
C655 a_36773_n5468 a_38403_n5503 0.213697f
C656 a_43892_n18820 a_44340_n18820 0.013276f
C657 a_42972_n20485 a_42884_n20388 0.285629f
C658 a_46020_n9032 a_46468_n9032 0.013276f
C659 a_43556_n10600 a_43196_n10644 0.087066f
C660 a_35849_n1192 a_35156_n325 0.016984f
C661 a_37372_n12212 a_37820_n12212 0.012882f
C662 a_28009_n12168 a_27639_n12537 0.374313f
C663 a_41764_n12168 a_41852_n12212 0.285629f
C664 a_40084_n10980 VDD 0.207208f
C665 a_46668_n14213 VDD 0.318039f
C666 a_37284_n15304 a_37732_n15304 0.013276f
C667 a_31292_n2804 a_30555_n2729 0.123873f
C668 a_24631_n3588 a_29856_n1121 0.035818f
C669 a_32468_n17252 VDD 0.216859f
C670 a_39076_n4328 a_39524_n4328 0.013276f
C671 a_40652_n1572 a_46243_769 0.033574f
C672 a_30372_376 a_30576_376 0.033243f
C673 a_46556_n20052 VDD 0.332067f
C674 a_43220_n5896 a_42860_n5940 0.087174f
C675 a_32220_n18484 a_32668_n18484 0.012882f
C676 a_36164_n18440 a_36252_n18484 0.285629f
C677 a_40956_n7508 CLK 0.010802f
C678 a_22948_n20008 a_22588_n20052 0.087066f
C679 a_22712_n7420 a_24233_n8684 0.019902f
C680 a_43420_n1669 VDD 0.330603f
C681 a_39164_n9076 a_39276_n9509 0.026339f
C682 a_42884_n20388 a_43332_n20388 0.013276f
C683 a_42996_n4708 VDD 0.208155f
C684 a_47004_n10644 a_47452_n10644 0.012222f
C685 a_46916_n12168 a_46556_n12212 0.086742f
C686 a_35268_n12168 VDD 0.127844f
C687 a_44004_n13736 a_44092_n13780 0.285629f
C688 a_21604_n708 a_21916_n1975 0.032513f
C689 a_40060_n13780 a_40508_n13780 0.012882f
C690 a_23360_n15233 VDD 0.826435f
C691 a_44452_n15304 a_44092_n15348 0.086635f
C692 a_39760_n4 VDD 0.01042f
C693 a_41092_n2760 a_41540_n2760 0.013276f
C694 a_27988_n20388 a_27085_n16132 0.042931f
C695 a_27988_n18440 VDD 0.203482f
C696 a_41852_n16916 a_42300_n16916 0.012882f
C697 a_28144_n4708 a_27190_n5112 0.010831f
C698 a_34012_n16916 a_33900_n17349 0.026339f
C699 a_38295_332 a_39056_820 0.042802f
C700 a_37947_332 a_38951_420 0.020455f
C701 a_45884_n20485 VDD 0.335211f
C702 a_47452_n5940 a_47900_n5940 0.012001f
C703 a_39524_n18440 a_39164_n18484 0.087066f
C704 a_29444_n20008 a_29892_n20008 0.013276f
C705 a_22220_n12996 a_25724_n14564 0.890094f
C706 a_38733_n5431 VDD 0.595386f
C707 a_29332_n11301 a_31544_n11296 0.042802f
C708 a_46668_n101 a_46580_n4 0.285629f
C709 a_46108_n9076 VDD 0.318654f
C710 a_27744_n12908 a_27639_n12537 0.536965f
C711 a_42748_n12212 a_42636_n12645 0.026339f
C712 a_26635_n12996 a_27535_n12493 0.116059f
C713 a_40508_n12212 VDD 0.315469f
C714 a_40420_n15304 VDD 0.205948f
C715 a_37859_377 a_41988_n2760 0.013991f
C716 a_35356_n18484 VDD 0.315469f
C717 a_22052_1944 a_25759_1944 0.034166f
C718 a_46243_769 a_46573_841 0.538085f
C719 a_46244_n20388 VDD 0.207333f
C720 a_35356_n18484 a_35244_n18917 0.026339f
C721 a_46020_n18440 a_46468_n18440 0.013276f
C722 a_30320_n6636 a_30808_n6334 0.08126f
C723 a_29559_n6456 a_30111_n6221 0.119687f
C724 a_36612_n20008 a_36252_n20052 0.086635f
C725 a_23564_n8292 a_21872_n9394 0.036893f
C726 a_22712_n7420 a_24965_n9860 0.047499f
C727 a_41740_n7941 a_42100_n7844 0.087066f
C728 a_44228_n2760 VDD 0.214978f
C729 a_24573_n9860 a_23816_n10112 0.032797f
C730 a_34392_n9815 a_28335_n10644 0.196648f
C731 a_42636_n14213 CLK 0.01698f
C732 a_22016_n6276 VDD 0.013678f
C733 a_41740_n11077 a_42188_n11077 0.012882f
C734 a_32581_n9860 VDD 0.49268f
C735 a_28492_n12548 VDD 0.298894f
C736 a_31789_n14564 a_32413_n14564 0.104193f
C737 a_45660_n13780 a_45772_n14213 0.026339f
C738 a_23954_n2020 a_24315_n2759 0.112057f
C739 a_26755_n16132 VDD 0.325638f
C740 a_21692_2431 a_29332_1243 0.183927f
C741 a_46108_n18484 VDD 0.318654f
C742 a_28972_n17349 a_28884_n17252 0.285629f
C743 a_39276_n17349 a_39724_n17349 0.012882f
C744 a_45212_n4372 a_45324_n4805 0.026339f
C745 a_42300_n18484 a_42188_n18917 0.026339f
C746 a_41740_n6373 a_41652_n6276 0.285629f
C747 a_46668_n6373 a_47116_n6373 0.012882f
C748 a_23479_n5156 a_26531_n8639 0.02172f
C749 a_43108_n20008 a_43556_n20008 0.013276f
C750 a_39524_n20008 a_39612_n20052 0.285629f
C751 a_42772_n4 VDD 0.207805f
C752 a_44004_n1192 VDD 1.30784f
C753 a_38292_n9412 a_38740_n9412 0.013276f
C754 a_46220_n9509 a_46132_n9412 0.285629f
C755 a_44876_n11077 a_44788_n10980 0.285629f
C756 a_28437_n13705 a_28040_n12493 0.026252f
C757 a_41652_n9412 VDD 0.205948f
C758 a_38604_n12645 a_38964_n12548 0.086905f
C759 a_25831_n12996 a_27302_n13160 0.020272f
C760 a_26635_n12996 a_26266_n13736 0.032175f
C761 a_26239_n12996 a_26470_n13736 0.013627f
C762 a_47564_n12645 a_48012_n12645 0.012882f
C763 a_34796_n14213 a_35156_n14116 0.087066f
C764 a_27988_n4328 a_31348_n1931 0.486192f
C765 a_33364_n15684 VDD 0.227717f
C766 a_47116_n15781 a_47564_n15781 0.012882f
C767 a_35800_n3456 a_36112_n3456 0.119687f
C768 a_38828_n15781 a_38740_n15684 0.285629f
C769 a_35568_n4 a_37680_n320 0.277491f
C770 a_41292_n18917 VDD 0.318502f
C771 a_22544_n4690 a_21604_n5412 0.012114f
C772 a_39724_n17349 a_40084_n17252 0.087066f
C773 a_22444_n5156 a_22264_n5852 0.054544f
C774 a_27988_n4328 a_21872_n9394 0.017768f
C775 a_24380_n18917 a_24740_n18820 0.087174f
C776 a_37932_n18917 a_38380_n18917 0.012882f
C777 a_38964_n7844 a_39076_n9032 0.026657f
C778 a_27485_n8500 a_21872_n9394 0.465551f
C779 a_39412_n3140 VDD 0.136232f
C780 a_22016_n10529 a_22364_n10512 0.401636f
C781 a_21604_n10116 a_22568_n10512 0.08126f
C782 a_37844_1564 VDD 1.00855f
C783 a_28335_n10644 a_32732_n10556 0.020277f
C784 a_47476_n10980 a_47924_n10980 0.013276f
C785 a_22500_n1976 a_28456_n364 0.133975f
C786 a_41988_n20388 CLK 0.014911f
C787 a_27302_n13160 VDD 0.574098f
C788 a_36948_n14116 a_37396_n14116 0.013276f
C789 a_45772_n14213 a_45684_n14116 0.285629f
C790 a_32860_n2020 a_32100_n1976 0.392453f
C791 a_22500_n1976 a_22568_n1104 0.021245f
C792 a_25544_n16412 VDD 0.528733f
C793 a_25600_n5895 a_26047_n4328 0.02863f
C794 a_45324_n3237 a_45772_n3237 0.012882f
C795 a_41292_n3237 a_41204_n3140 0.285629f
C796 a_35064_1506 a_35324_1564 0.66083f
C797 a_36052_n18820 VDD 0.206648f
C798 a_34576_1204 a_37396_1205 0.045724f
C799 a_45772_n4805 a_45684_n4708 0.285629f
C800 a_40084_n17252 a_40532_n17252 0.013276f
C801 a_30396_n7508 a_30036_n7464 0.582861f
C802 a_35692_n18917 a_35604_n18820 0.285629f
C803 a_31100_n20485 a_31548_n20485 0.013103f
C804 a_44540_n20052 a_44540_n20485 0.05841f
C805 a_25831_n11428 a_25880_n11708 0.01241f
C806 a_44540_n7508 VDD 0.353322f
C807 a_27281_n16854 a_27804_n14165 0.01857f
C808 a_25573_n12167 a_25160_n14816 0.015136f
C809 a_42300_n10644 VDD 0.315469f
C810 a_39972_n13736 VDD 0.207563f
C811 a_45660_n1669 a_45572_n1572 0.285629f
C812 a_41764_n16872 VDD 0.206217f
C813 a_22948_n16872 a_23036_n16916 0.285629f
C814 a_24631_n3588 a_22052_n4708 0.012444f
C815 a_37859_377 a_39056_820 0.038103f
C816 a_21692_n20052 VDD 0.317437f
C817 a_34708_n17252 a_34820_n18440 0.026657f
C818 a_21604_n5412 a_22016_n5825 0.536965f
C819 a_46220_n18917 a_46580_n18820 0.087066f
C820 a_38733_n727 VDD 0.599022f
C821 a_39524_n9032 a_39164_n9076 0.087066f
C822 a_31548_n20485 a_31460_n20388 0.285629f
C823 a_43108_n9032 a_43556_n9032 0.013276f
C824 a_44540_n4372 VDD 0.353742f
C825 a_22264_n8988 a_21872_n12530 0.021426f
C826 a_24965_n9860 a_23212_n12124 0.039052f
C827 a_25020_n11383 a_31544_n11296 0.022355f
C828 a_32581_n9860 a_32158_n12212 0.024011f
C829 a_39352_464 VDD 0.245198f
C830 a_40396_n7941 VDD 0.333825f
C831 a_47924_n10980 a_47812_n12168 0.026657f
C832 a_31961_n11340 VDD 0.465287f
C833 a_44340_n12548 a_44452_n13736 0.026657f
C834 a_30555_n13780 a_31664_n13292 0.019043f
C835 a_42548_n14116 a_42660_n15304 0.026657f
C836 a_37221_n3543 a_39357_n2228 0.522698f
C837 a_35849_n1192 a_34895_n1192 0.019369f
C838 a_31212_n17349 VDD 0.336066f
C839 a_31684_n16872 a_31324_n16916 0.087174f
C840 a_35356_n20052 VDD 0.296789f
C841 a_35849_n1192 a_30104_n1148 0.034422f
C842 a_41652_n17252 a_41764_n18440 0.026657f
C843 a_36773_n5468 a_37732_n5896 0.021708f
C844 a_45236_n4708 a_45124_n5896 0.026657f
C845 a_41404_n7508 a_41852_n7508 0.012882f
C846 a_31460_n20388 a_31908_n20388 0.013276f
C847 a_42524_n20485 a_42884_n20388 0.087174f
C848 a_43108_n10600 a_43196_n10644 0.285629f
C849 a_39164_n10644 a_39612_n10644 0.012882f
C850 a_41764_n12168 a_41404_n12212 0.087066f
C851 a_39636_n10980 VDD 0.210107f
C852 a_36588_n13780 a_37284_n13736 0.012267f
C853 a_46220_n14213 VDD 0.31977f
C854 a_32020_n17252 VDD 0.213721f
C855 a_38628_n16872 a_39076_n16872 0.013276f
C856 a_34271_376 a_31076_376 0.020162f
C857 a_40652_n1572 a_45572_376 0.081681f
C858 a_46108_n20052 VDD 0.333671f
C859 a_42772_n5896 a_42860_n5940 0.285629f
C860 a_36164_n18440 a_35804_n18484 0.087066f
C861 a_39612_n7508 a_39500_n7941 0.026339f
C862 a_26084_n20008 a_26532_n20008 0.013276f
C863 a_22500_n20008 a_22588_n20052 0.285629f
C864 a_36500_n18820 a_36612_n20008 0.026657f
C865 a_42244_n1572 VDD 0.594443f
C866 a_25831_n11428 a_25020_n11383 0.088363f
C867 a_42548_n4708 VDD 0.208155f
C868 a_21772_n9860 a_21872_n12530 1.17793f
C869 a_35804_n12212 a_35916_n12645 0.026339f
C870 a_46468_n12168 a_46556_n12212 0.285629f
C871 a_33910_n12146 VDD 0.317492f
C872 a_44004_n13736 a_43644_n13780 0.087066f
C873 a_22140_n15348 VDD 0.30145f
C874 a_40060_n15348 a_40508_n15348 0.012882f
C875 a_23507_n2759 a_25759_n3544 0.04701f
C876 a_44004_n15304 a_44092_n15348 0.285629f
C877 a_22164_n2760 a_27932_n3543 0.198038f
C878 a_27540_n18440 VDD 0.209136f
C879 a_41404_n4372 a_41852_n4372 0.013103f
C880 a_37947_332 a_39056_820 0.019043f
C881 a_45436_n20485 VDD 0.337745f
C882 a_42660_n18440 a_43108_n18440 0.013276f
C883 a_39076_n18440 a_39164_n18484 0.285629f
C884 a_43444_n18820 a_43556_n20008 0.026657f
C885 a_37260_n7941 a_37708_n7941 0.013103f
C886 a_25547_n2445 VDD 1.03982f
C887 a_38403_n5503 VDD 0.349684f
C888 a_46220_n101 a_46580_n4 0.086905f
C889 a_45660_n9076 VDD 0.320877f
C890 a_26983_n12728 a_27639_n12537 0.510371f
C891 a_40060_n12212 VDD 0.316003f
C892 a_47452_n13780 a_47900_n13780 0.012001f
C893 a_39972_n15304 VDD 0.207295f
C894 a_34232_n2272 a_33588_n3461 0.035006f
C895 a_38268_n15348 a_38380_n15781 0.026339f
C896 a_32860_n2020 a_32911_n4240 0.050051f
C897 a_34908_n18484 VDD 0.315469f
C898 a_40508_n16916 a_40620_n17349 0.026339f
C899 a_28076_n17349 a_28524_n17349 0.013103f
C900 a_22444_n5156 a_22544_n4690 0.026393f
C901 a_45796_n20388 VDD 0.209377f
C902 a_29211_n6724 a_30111_n6221 0.116059f
C903 a_30320_n6636 a_30215_n6265 0.536965f
C904 a_47004_n5940 a_47116_n6373 0.026339f
C905 a_36164_n20008 a_36252_n20052 0.285629f
C906 a_32220_n20052 a_32668_n20052 0.012882f
C907 a_41740_n7941 a_41652_n7844 0.285629f
C908 a_43780_n2760 VDD 0.20719f
C909 a_33494_n9860 a_28335_n10644 0.18058f
C910 a_42636_n9509 a_43084_n9509 0.012882f
C911 a_42188_n14213 CLK 0.047331f
C912 a_31961_n11340 a_32158_n12212 0.151669f
C913 a_32189_n9860 VDD 0.748313f
C914 a_36364_n12645 a_36812_n12645 0.013103f
C915 a_28040_n12493 VDD 0.244473f
C916 a_28752_n15348 a_32413_n14564 0.464356f
C917 a_23954_n2020 a_24578_n2020 0.107109f
C918 a_23542_n1754 a_24315_n2759 0.013135f
C919 a_33077_n1191 a_36388_n1572 0.038799f
C920 a_24752_n16132 VDD 0.577675f
C921 a_22164_n2760 a_27540_n3797 0.014746f
C922 a_47452_n15348 a_47564_n15781 0.026339f
C923 a_36140_n15781 a_36588_n15781 0.012882f
C924 a_45660_n18484 VDD 0.320877f
C925 a_28524_n17349 a_28884_n17252 0.087174f
C926 a_26956_n18917 a_27404_n18917 0.012882f
C927 a_41292_n6373 a_41652_n6276 0.087066f
C928 a_22444_n5156 a_21872_n9394 0.011031f
C929 a_39524_n20008 a_39164_n20052 0.087066f
C930 a_45236_n7844 a_45684_n7844 0.013276f
C931 a_27337_n3140 VDD 0.405299f
C932 a_45772_n9509 a_46132_n9412 0.087066f
C933 a_29992_n11150 a_28927_n10160 0.023082f
C934 a_39412_n6276 VDD 0.130441f
C935 a_44428_n11077 a_44788_n10980 0.087066f
C936 a_41204_n9412 VDD 0.226701f
C937 a_26239_n12996 a_26266_n13736 0.013163f
C938 a_23564_n11428 a_25472_n14816 0.038162f
C939 a_38604_n12645 a_38516_n12548 0.285629f
C940 a_24684_n16432 a_23608_n15260 0.085501f
C941 a_34796_n14213 a_34708_n14116 0.285629f
C942 a_43084_n14213 a_43532_n14213 0.012882f
C943 a_45660_n1236 a_45660_n1669 0.05841f
C944 a_23564_n17700 VDD 1.5551f
C945 a_38380_n15781 a_38740_n15684 0.087066f
C946 a_35800_n3456 a_36217_n3500 0.633318f
C947 a_35568_n4 a_37785_n364 0.020455f
C948 a_40620_n18917 VDD 0.343849f
C949 a_27988_n4328 a_27485_n8500 0.013804f
C950 a_47564_n101 a_47476_n4 0.285629f
C951 a_39724_n17349 a_39636_n17252 0.285629f
C952 a_28884_n17252 a_29332_n17252 0.013276f
C953 OUT[1] OUT[2] 0.0571f
C954 a_22444_n5156 a_22016_n5825 0.0169f
C955 VDD OUT[3] 1.32407f
C956 a_24380_n18917 a_24292_n18820 0.285629f
C957 a_46580_n6276 a_47028_n6276 0.013276f
C958 a_23816_n8544 a_24128_n8544 0.119687f
C959 a_46020_n20008 a_46468_n20008 0.013276f
C960 a_26861_n8567 a_21872_n9394 0.079265f
C961 a_48012_n3237 VDD 0.343887f
C962 a_24965_n9860 a_23564_n11428 0.073631f
C963 a_28335_n10644 a_31872_n10529 0.040035f
C964 a_22016_n10529 a_22876_n10556 0.882105f
C965 a_21604_n10116 a_22364_n10512 0.011851f
C966 a_37396_1205 VDD 0.477937f
C967 a_35156_n325 a_35568_n4 0.536965f
C968 a_31799_n7508 VDD 1.34931f
C969 a_30808_n10116 VDD 0.299659f
C970 a_26470_n13736 VDD 0.736231f
C971 a_45324_n14213 a_45684_n14116 0.087066f
C972 a_32636_n2020 a_32100_n1976 0.44798f
C973 a_23932_n16916 VDD 0.324594f
C974 a_25600_n5895 a_25423_n4328 0.073975f
C975 a_35064_1506 a_34872_1619 0.934191f
C976 a_35604_n18820 VDD 0.206648f
C977 a_45324_n4805 a_45684_n4708 0.087066f
C978 a_39076_n4708 a_39524_n4708 0.013276f
C979 a_42548_n6276 a_42660_n7464 0.026657f
C980 a_25972_n6276 a_27597_n8292 0.056553f
C981 a_21604_n18820 a_22052_n18820 0.013276f
C982 a_29476_n6980 a_30036_n7464 0.302602f
C983 a_35244_n18917 a_35604_n18820 0.087066f
C984 a_45684_n7844 a_45572_n9032 0.026657f
C985 a_28435_n10599 a_29444_n10116 0.011241f
C986 a_29992_n11150 a_29332_n11301 0.104374f
C987 a_28927_n10160 a_28247_n10599 0.163112f
C988 a_42548_n9412 a_42660_n10600 0.026657f
C989 a_44092_n7508 VDD 0.3211f
C990 a_27281_n16854 a_27192_n14286 0.390977f
C991 a_25573_n12167 a_25577_n14956 0.012803f
C992 a_41204_n10980 a_41316_n12168 0.026657f
C993 a_41852_n10644 VDD 0.315469f
C994 a_41864_1394 a_42948_n1976 0.051432f
C995 a_39524_n13736 VDD 0.209768f
C996 a_45212_n1669 a_45572_n1572 0.087174f
C997 a_47476_n14116 a_47924_n14116 0.013276f
C998 a_34708_n14116 a_34708_n15304 0.05841f
C999 a_27988_n4328 a_27628_n3841 0.054396f
C1000 a_41316_n16872 VDD 0.206217f
C1001 a_22948_n16872 a_22588_n16916 0.086905f
C1002 a_47028_n3140 a_47476_n3140 0.013276f
C1003 a_28772_n20008 VDD 0.213111f
C1004 a_24492_n5156 a_25972_n6276 0.535858f
C1005 a_23844_n18440 a_24292_n18440 0.013276f
C1006 a_22220_n9860 a_21812_n6643 0.280456f
C1007 a_46220_n18917 a_46132_n18820 0.285629f
C1008 a_38180_n7464 a_38628_n7464 0.013276f
C1009 a_38403_n799 VDD 0.351691f
C1010 a_42076_n20485 a_42524_n20485 0.013103f
C1011 a_39076_n9032 a_39164_n9076 0.285629f
C1012 a_31100_n20485 a_31460_n20388 0.087174f
C1013 a_23564_n8292 a_22016_n10529 0.027741f
C1014 a_44092_n4372 VDD 0.32119f
C1015 a_34652_n11391 a_33900_n11428 0.059328f
C1016 a_39948_n7941 VDD 0.315604f
C1017 a_31544_n11296 VDD 1.34308f
C1018 a_37221_n3543 a_38733_n2295 0.092164f
C1019 a_22820_n2804 a_23507_n2759 0.05696f
C1020 a_30764_n17349 VDD 0.321135f
C1021 a_34372_n16872 a_34820_n16872 0.013276f
C1022 a_31236_n16872 a_31324_n16916 0.285629f
C1023 a_42996_n3140 a_43108_n4328 0.026657f
C1024 a_34908_n20052 VDD 0.296789f
C1025 a_36773_n5468 a_37284_n5896 0.019585f
C1026 a_43444_n18820 a_43892_n18820 0.013276f
C1027 a_45572_n9032 a_46020_n9032 0.013276f
C1028 a_42524_n20485 a_42436_n20388 0.285629f
C1029 a_32132_n4708 VDD 0.650715f
C1030 a_28927_n10160 a_30296_n10980 0.039602f
C1031 a_43108_n10600 a_42748_n10644 0.087066f
C1032 a_47924_n7844 VDD 0.21239f
C1033 a_41316_n12168 a_41404_n12212 0.285629f
C1034 a_39188_n10980 VDD 0.211835f
C1035 a_26431_n1192 a_25524_n708 0.019505f
C1036 a_45772_n14213 VDD 0.321879f
C1037 a_36588_n15348 a_37284_n15304 0.012267f
C1038 a_31572_n17252 VDD 0.237441f
C1039 a_40652_n1572 a_45124_376 0.014911f
C1040 a_45660_n20052 VDD 0.335894f
C1041 a_28492_332 a_30104_n1148 0.963309f
C1042 a_42772_n5896 a_42412_n5940 0.087174f
C1043 a_35716_n18440 a_35804_n18484 0.285629f
C1044 a_31772_n18484 a_32220_n18484 0.012882f
C1045 a_22500_n20008 a_22140_n20052 0.087066f
C1046 a_41684_n1976 VDD 0.556603f
C1047 a_42436_n20388 a_42884_n20388 0.013276f
C1048 a_38716_n9076 a_38828_n9509 0.026339f
C1049 a_42100_n4708 VDD 0.208155f
C1050 a_21772_n9860 a_23619_n12996 0.012648f
C1051 a_46556_n10644 a_47004_n10644 0.012222f
C1052 a_25831_n11428 VDD 1.22327f
C1053 a_46468_n12168 a_46108_n12212 0.086905f
C1054 a_33686_n11592 VDD 0.592071f
C1055 a_39612_n13780 a_40060_n13780 0.012882f
C1056 a_27820_n16432 a_28752_n15348 0.068955f
C1057 a_34895_n1192 a_33077_n1191 0.012001f
C1058 a_43556_n13736 a_43644_n13780 0.285629f
C1059 a_21692_n15348 VDD 0.300735f
C1060 a_44004_n15304 a_43644_n15348 0.087066f
C1061 a_40644_n2760 a_41092_n2760 0.013276f
C1062 a_23507_n2759 a_25237_n4327 0.040355f
C1063 a_27092_n18440 VDD 0.131804f
C1064 a_41404_n16916 a_41852_n16916 0.012882f
C1065 a_33564_n16916 a_33452_n17349 0.026339f
C1066 a_44988_n20485 VDD 0.372934f
C1067 a_39076_n18440 a_38716_n18484 0.087066f
C1068 a_47004_n5940 a_47452_n5940 0.012222f
C1069 a_22444_n5156 a_23564_n8292 0.012889f
C1070 a_28860_n20052 a_29444_n20008 0.016748f
C1071 a_24771_n2804 VDD 0.320099f
C1072 a_47900_n9076 a_48012_n9509 0.026339f
C1073 a_42604_n2020 a_45684_n4 0.014194f
C1074 a_37732_n5896 VDD 0.212864f
C1075 a_29332_n11301 a_30296_n10980 0.08126f
C1076 a_45212_n9076 VDD 0.342281f
C1077 a_42300_n12212 a_42188_n12645 0.026339f
C1078 a_26635_n12996 a_27639_n12537 0.020455f
C1079 a_39612_n12212 VDD 0.31906f
C1080 a_42972_n1236 a_43556_n661 0.04398f
C1081 a_39524_n15304 VDD 0.209499f
C1082 a_34649_n2412 a_33588_n3461 0.080901f
C1083 a_47452_n15348 a_47900_n15348 0.012001f
C1084 a_34460_n18484 VDD 0.315469f
C1085 a_45348_n20388 VDD 0.213014f
C1086 a_45572_n18440 a_46020_n18440 0.013276f
C1087 a_34908_n18484 a_34796_n18917 0.026339f
C1088 a_29559_n6456 a_30215_n6265 0.510371f
C1089 a_41292_n7941 a_41652_n7844 0.087066f
C1090 a_36164_n20008 a_35804_n20052 0.087066f
C1091 a_43332_n2760 VDD 0.205276f
C1092 a_32581_n9860 a_28335_n10644 0.033343f
C1093 a_29992_n11150 a_25020_n11383 0.210577f
C1094 a_23619_n6724 VDD 0.309736f
C1095 a_41292_n11077 a_41740_n11077 0.012882f
C1096 a_31544_n11296 a_32158_n12212 0.019626f
C1097 a_31565_n9860 VDD 0.618081f
C1098 a_27535_n12493 VDD 0.022335f
C1099 a_28752_n15348 a_31789_n14564 0.081658f
C1100 a_45212_n13780 a_45324_n14213 0.026339f
C1101 a_24088_n16087 VDD 0.449834f
C1102 a_27988_n4328 a_22444_n5156 0.047648f
C1103 a_26383_n2968 a_26607_n3544 0.538085f
C1104 a_22164_n2760 a_28144_n4708 0.428203f
C1105 a_28736_1944 a_28583_n3140 0.037814f
C1106 a_21692_2431 a_28153_1204 0.17465f
C1107 a_37859_377 a_39748_2475 0.518272f
C1108 a_45212_n18484 VDD 0.342281f
C1109 a_28524_n17349 a_28436_n17252 0.285629f
C1110 a_38828_n17349 a_39276_n17349 0.012882f
C1111 a_41852_n18484 a_41740_n18917 0.026339f
C1112 a_46220_n6373 a_46668_n6373 0.012882f
C1113 a_41292_n6373 a_41204_n6276 0.285629f
C1114 a_39076_n20008 a_39164_n20052 0.285629f
C1115 a_42660_n20008 a_43108_n20008 0.013276f
C1116 a_45772_n9509 a_45684_n9412 0.285629f
C1117 a_37844_n9412 a_38292_n9412 0.013276f
C1118 a_44428_n11077 a_44340_n10980 0.285629f
C1119 a_36500_n10980 a_36948_n10980 0.013276f
C1120 a_28437_n13705 a_28232_n12606 0.01568f
C1121 a_40532_n9412 VDD 0.212412f
C1122 a_25831_n12996 a_26266_n13736 0.018815f
C1123 a_38156_n12645 a_38516_n12548 0.086905f
C1124 a_47116_n12645 a_47564_n12645 0.012882f
C1125 a_26239_n12996 a_25642_n13736 0.023071f
C1126 a_30584_n1954 a_31348_n1931 0.238627f
C1127 a_34348_n14213 a_34708_n14116 0.087066f
C1128 a_38380_n15781 a_38292_n15684 0.285629f
C1129 a_46668_n15781 a_47116_n15781 0.012882f
C1130 a_35568_n4 a_37368_n320 0.510371f
C1131 a_36428_n53 a_36324_n4 0.026665f
C1132 a_40172_n18917 VDD 0.315469f
C1133 a_22444_n5156 a_21604_n5412 0.047699f
C1134 a_39276_n17349 a_39636_n17252 0.087066f
C1135 a_40060_n4805 a_40508_n4805 0.012222f
C1136 a_47116_n101 a_47476_n4 0.086742f
C1137 a_37484_n18917 a_37932_n18917 0.012882f
C1138 a_23932_n18917 a_24292_n18820 0.087174f
C1139 a_24233_n8684 a_24128_n8544 0.116059f
C1140 a_26531_n8639 a_21872_n9394 0.02976f
C1141 a_26861_n8567 a_27485_n8500 0.104193f
C1142 a_38516_n7844 a_38628_n9032 0.026657f
C1143 a_47564_n3237 VDD 0.315945f
C1144 a_21604_n10116 a_22876_n10556 0.05539f
C1145 a_31451_n7508 VDD 0.517973f
C1146 a_47028_n10980 a_47476_n10980 0.013276f
C1147 a_26266_n13736 VDD 0.593638f
C1148 a_27192_n14286 a_27988_n20388 0.121786f
C1149 a_45324_n14213 a_45236_n14116 0.285629f
C1150 a_36500_n14116 a_36948_n14116 0.013276f
C1151 a_22500_n1976 a_22876_n1148 0.062137f
C1152 a_23484_n16916 VDD 0.317396f
C1153 a_40396_n3237 a_40308_n3140 0.285629f
C1154 a_44876_n3237 a_45324_n3237 0.012882f
C1155 a_34471_1575 a_34872_1619 0.882105f
C1156 a_35156_n18820 VDD 0.206648f
C1157 a_34576_1204 a_35849_n1192 0.11373f
C1158 a_39636_n17252 a_40084_n17252 0.013276f
C1159 a_45324_n4805 a_45236_n4708 0.285629f
C1160 a_35244_n18917 a_35156_n18820 0.285629f
C1161 a_29476_n6980 a_30396_n7508 0.0144f
C1162 a_25972_n6276 a_26973_n8292 0.022851f
C1163 a_30652_n20485 a_31100_n20485 0.013103f
C1164 a_28437_n13705 a_28247_n10599 0.124155f
C1165 a_43644_n7508 VDD 0.319164f
C1166 a_27281_n16854 a_26944_n14116 0.034477f
C1167 a_41404_n10644 VDD 0.315469f
C1168 a_39076_n13736 VDD 0.211682f
C1169 a_45212_n1669 a_45124_n1572 0.285629f
C1170 a_40868_n16872 VDD 0.208618f
C1171 a_22500_n16872 a_22588_n16916 0.285629f
C1172 a_37859_377 a_38295_332 0.034316f
C1173 a_28324_n20008 VDD 0.206367f
C1174 a_22444_n5156 a_29123_n6679 0.024586f
C1175 a_23887_n5156 a_25972_n6276 0.088523f
C1176 a_34260_n17252 a_34372_n18440 0.026657f
C1177 a_45772_n18917 a_46132_n18820 0.087066f
C1178 a_32244_n18820 a_32692_n18820 0.013276f
C1179 a_26861_n8567 a_26470_n9322 0.018566f
C1180 a_42660_n9032 a_43108_n9032 0.013276f
C1181 a_25573_n12167 a_21772_n9860 0.019142f
C1182 a_39076_n9032 a_38716_n9076 0.087066f
C1183 a_31100_n20485 a_31012_n20388 0.285629f
C1184 a_39556_n4 VDD 0.591706f
C1185 a_43644_n4372 VDD 0.319254f
C1186 a_24965_n9860 a_22352_n12097 0.035943f
C1187 a_25020_n11383 a_30296_n10980 0.026694f
C1188 a_38847_464 VDD 0.024358f
C1189 a_39500_n7941 VDD 0.317865f
C1190 a_47476_n10980 a_47364_n12168 0.026657f
C1191 a_30500_n10980 VDD 0.298894f
C1192 a_30555_n13780 a_30903_n13780 0.633318f
C1193 a_43892_n12548 a_44004_n13736 0.026657f
C1194 a_26532_n14437 VDD 1.7995f
C1195 a_42100_n14116 a_42212_n15304 0.026657f
C1196 a_37221_n3543 a_38403_n2367 0.013216f
C1197 a_30316_n17349 VDD 0.318699f
C1198 a_31236_n16872 a_30876_n16916 0.087174f
C1199 a_34460_n20052 VDD 0.296789f
C1200 a_36773_n5468 a_29612_n8292 0.4072f
C1201 a_41204_n17252 a_41316_n18440 0.026657f
C1202 a_28076_n18484 a_28524_n18484 0.012552f
C1203 a_40956_n7508 a_41404_n7508 0.012882f
C1204 a_42076_n20485 a_42436_n20388 0.087174f
C1205 a_25831_n11428 a_31235_n9860 0.016809f
C1206 a_31919_n9032 a_32189_n9860 0.025177f
C1207 a_31012_n20388 a_31460_n20388 0.013276f
C1208 a_42660_n10600 a_42748_n10644 0.285629f
C1209 a_38716_n10644 a_39164_n10644 0.012882f
C1210 a_47476_n7844 VDD 0.206217f
C1211 a_41316_n12168 a_40956_n12212 0.087066f
C1212 a_38740_n10980 VDD 0.214497f
C1213 a_24684_n16432 a_25544_n16412 0.015911f
C1214 a_36140_n13780 a_36588_n13780 0.012001f
C1215 a_45324_n14213 VDD 0.324845f
C1216 a_31124_n17252 VDD 0.216838f
C1217 a_38180_n16872 a_38628_n16872 0.013276f
C1218 a_33533_908 a_31076_376 0.024415f
C1219 a_45212_n20052 VDD 0.358183f
C1220 a_42324_n5896 a_42412_n5940 0.285629f
C1221 a_35716_n18440 a_35356_n18484 0.087066f
C1222 a_25636_n20008 a_26084_n20008 0.013276f
C1223 a_22052_n20008 a_22140_n20052 0.285629f
C1224 a_36052_n18820 a_36164_n20008 0.026657f
C1225 a_39164_n7508 a_39052_n7941 0.026339f
C1226 a_22712_n7420 a_22568_n8944 0.060288f
C1227 a_41292_n1669 VDD 0.331215f
C1228 a_26266_n9240 a_26470_n9322 0.499501f
C1229 a_41652_n4708 VDD 0.208155f
C1230 a_28435_n10599 a_33364_n11384 0.523618f
C1231 a_21772_n9860 a_21772_n12996 0.052109f
C1232 a_34092_n9076 VDD 0.490675f
C1233 a_46020_n12168 a_46108_n12212 0.285629f
C1234 a_47364_n12168 a_47812_n12168 0.013276f
C1235 a_35356_n12212 a_35468_n12645 0.026339f
C1236 a_32854_n12168 VDD 0.768417f
C1237 a_41864_1394 a_43555_n452 0.211511f
C1238 a_43556_n13736 a_43196_n13780 0.087066f
C1239 a_34271_n1192 a_33077_n1191 0.015807f
C1240 a_22948_n14820 VDD 1.88874f
C1241 a_39612_n15348 a_40060_n15348 0.012882f
C1242 a_43556_n15304 a_43644_n15348 0.285629f
C1243 a_26084_n18440 VDD 0.213959f
C1244 a_40956_n4372 a_41404_n4372 0.013103f
C1245 a_47028_n4 a_47476_n4 0.013276f
C1246 a_37947_332 a_38295_332 0.633318f
C1247 a_44540_n20485 VDD 0.309901f
C1248 a_38628_n18440 a_38716_n18484 0.285629f
C1249 a_42212_n18440 a_42660_n18440 0.013276f
C1250 a_36812_n7941 a_37260_n7941 0.013103f
C1251 a_42996_n18820 a_43108_n20008 0.026657f
C1252 a_31235_n9860 a_31565_n9860 0.538085f
C1253 a_37284_n5896 VDD 0.22875f
C1254 a_29332_n11301 a_30092_n10980 0.011851f
C1255 a_47812_n9032 VDD 0.211703f
C1256 a_39164_n12212 VDD 0.320885f
C1257 a_47004_n13780 a_47452_n13780 0.012222f
C1258 a_39076_n15304 VDD 0.211414f
C1259 a_32860_n2020 a_33015_n4284 0.024538f
C1260 a_43868_n2804 a_44316_n2804 0.012001f
C1261 a_37820_n15348 a_37932_n15781 0.026339f
C1262 a_34012_n18484 VDD 0.315469f
C1263 a_21604_2475 a_22052_1944 0.195233f
C1264 a_40060_n16916 a_40172_n17349 0.026339f
C1265 a_44900_n20388 VDD 0.231097f
C1266 a_46556_n5940 a_46668_n6373 0.026339f
C1267 a_29211_n6724 a_30215_n6265 0.020455f
C1268 a_41292_n7941 a_41204_n7844 0.285629f
C1269 a_24752_n8292 a_23816_n8544 0.034291f
C1270 a_31772_n20052 a_32220_n20052 0.012882f
C1271 a_35716_n20008 a_35804_n20052 0.285629f
C1272 a_22712_n7420 a_22264_n10556 0.02716f
C1273 a_42884_n2760 VDD 0.203482f
C1274 a_42188_n9509 a_42636_n9509 0.012882f
C1275 a_25724_n14564 a_25020_n11383 0.032145f
C1276 a_22968_n6679 VDD 0.443295f
C1277 a_29992_n11150 VDD 0.563237f
C1278 a_35916_n12645 a_36364_n12645 0.013103f
C1279 a_28232_n12606 VDD 0.360568f
C1280 a_33077_n1191 a_35940_n1931 0.522468f
C1281 a_23542_n1754 a_23954_n2020 0.499501f
C1282 a_23036_n15781 VDD 0.337685f
C1283 a_25237_n4327 a_27932_n3543 0.044398f
C1284 a_47004_n15348 a_47116_n15781 0.026339f
C1285 a_35692_n15781 a_36140_n15781 0.012882f
C1286 a_21692_2431 a_27736_1248 0.035205f
C1287 a_47812_n18440 VDD 0.211703f
C1288 a_28076_n17349 a_28436_n17252 0.087174f
C1289 a_26508_n18917 a_26956_n18917 0.012882f
C1290 a_44788_n7844 a_45236_n7844 0.013276f
C1291 a_39076_n20008 a_38716_n20052 0.087066f
C1292 a_45324_n9509 a_45684_n9412 0.087066f
C1293 a_31936_n6592 VDD 0.012699f
C1294 a_43980_n11077 a_44340_n10980 0.087066f
C1295 a_28437_n13705 a_27639_n12537 0.018187f
C1296 a_28121_n10980 a_28009_n12168 0.716733f
C1297 a_40084_n9412 VDD 0.206509f
C1298 a_38156_n12645 a_38068_n12548 0.285629f
C1299 a_25831_n12996 a_25642_n13736 0.054625f
C1300 a_26563_n12212 a_26944_n14116 0.028187f
C1301 a_42636_n14213 a_43084_n14213 0.012882f
C1302 a_45212_n1236 a_45212_n1669 0.05841f
C1303 a_34348_n14213 a_34260_n14116 0.285629f
C1304 a_37932_n15781 a_38292_n15684 0.087066f
C1305 a_29560_n3544 a_31676_n3544 0.012389f
C1306 a_26488_1564 a_26692_1564 0.66083f
C1307 a_39724_n18917 VDD 0.318714f
C1308 a_39276_n17349 a_39188_n17252 0.285629f
C1309 a_28436_n17252 a_28884_n17252 0.013276f
C1310 a_36773_n5468 CLK 0.027619f
C1311 a_23932_n18917 a_23844_n18820 0.285629f
C1312 a_46132_n6276 a_46580_n6276 0.013276f
C1313 a_45572_n20008 a_46020_n20008 0.013276f
C1314 a_23816_n8544 a_21872_n9394 0.011035f
C1315 a_47116_n3237 VDD 0.315945f
C1316 a_21604_n10116 a_22016_n10529 0.536965f
C1317 a_21772_n9860 a_26547_n12951 0.030441f
C1318 a_35849_n1192 VDD 0.505017f
C1319 a_28335_n10644 a_30808_n10116 0.143614f
C1320 a_32158_n12212 a_32854_n12168 0.012508f
C1321 a_28247_n10599 VDD 0.976715f
C1322 a_33488_n12996 a_31664_n13292 0.035264f
C1323 a_39860_n12548 a_40308_n12548 0.013276f
C1324 a_25642_n13736 VDD 0.700645f
C1325 a_44876_n14213 a_45236_n14116 0.087066f
C1326 a_23036_n16916 VDD 0.315221f
C1327 a_25237_n4327 a_27540_n3797 0.010544f
C1328 a_40084_n15684 a_40532_n15684 0.013276f
C1329 a_39948_n3237 a_40308_n3140 0.086635f
C1330 a_34471_1575 a_34367_1619 0.277491f
C1331 a_34708_n18820 VDD 0.206648f
C1332 a_44876_n4805 a_45236_n4708 0.087066f
C1333 a_38628_n4708 a_39076_n4708 0.013276f
C1334 a_34796_n18917 a_35156_n18820 0.087066f
C1335 a_42100_n6276 a_42212_n7464 0.026657f
C1336 a_45236_n7844 a_45124_n9032 0.026657f
C1337 a_42100_n9412 a_42212_n10600 0.026657f
C1338 a_28132_376 VDD 0.607515f
C1339 a_43196_n7508 VDD 0.316157f
C1340 a_28121_n10980 a_27744_n12908 0.069119f
C1341 a_41864_1394 a_43885_n452 0.014413f
C1342 a_40956_n10644 VDD 0.330158f
C1343 a_22876_n13692 a_23816_n13248 0.056721f
C1344 a_38628_n13736 VDD 0.214632f
C1345 a_34260_n14116 a_34260_n15304 0.05841f
C1346 a_47028_n14116 a_47476_n14116 0.013276f
C1347 a_27988_n4328 a_31292_n2804 0.083325f
C1348 a_44764_n1669 a_45124_n1572 0.087174f
C1349 a_40420_n16872 VDD 0.205948f
C1350 a_46580_n3140 a_47028_n3140 0.013276f
C1351 a_22500_n16872 a_22140_n16916 0.086905f
C1352 a_41864_1394 a_43644_n705 0.066219f
C1353 a_37859_377 a_37947_332 0.134996f
C1354 a_43833_1204 a_43728_1248 0.116059f
C1355 a_27876_n20008 VDD 0.206367f
C1356 a_23479_n5156 a_25972_n6276 0.089753f
C1357 a_23396_n18440 a_23844_n18440 0.013276f
C1358 a_25972_n6276 a_29532_n10311 0.788503f
C1359 a_45772_n18917 a_45684_n18820 0.285629f
C1360 a_37732_n7464 a_38180_n7464 0.013276f
C1361 a_30652_n20485 a_31012_n20388 0.087174f
C1362 a_38628_n9032 a_38716_n9076 0.285629f
C1363 a_41628_n20485 a_42076_n20485 0.013103f
C1364 a_38996_n408 VDD 0.488533f
C1365 a_43196_n4372 VDD 0.316247f
C1366 a_39544_420 VDD 0.362151f
C1367 a_39052_n7941 VDD 0.32028f
C1368 a_32132_2428 OUT[1] 0.011446f
C1369 a_30296_n10980 VDD 0.364257f
C1370 a_24516_n14475 VDD 0.550044f
C1371 a_34248_n3310 a_32020_n2276 0.011844f
C1372 a_29868_n17349 VDD 0.330483f
C1373 a_42548_n3140 a_42660_n4328 0.026657f
C1374 a_33924_n16872 a_34372_n16872 0.013276f
C1375 a_30788_n16872 a_30876_n16916 0.285629f
C1376 a_35156_n325 a_36120_n4 0.08126f
C1377 a_34012_n20052 VDD 0.296789f
C1378 a_23404_816 a_23004_n2332 0.029237f
C1379 a_42996_n18820 a_43444_n18820 0.013276f
C1380 a_42076_n20485 a_41988_n20388 0.285629f
C1381 a_25831_n11428 a_30472_n9815 0.016163f
C1382 a_45124_n9032 a_45572_n9032 0.013276f
C1383 a_30136_n10600 a_29332_n11301 0.032782f
C1384 a_42660_n10600 a_42300_n10644 0.087066f
C1385 a_33508_n408 a_34068_n4 0.302602f
C1386 a_47028_n7844 VDD 0.206217f
C1387 a_29540_n11728 a_27744_n12908 0.029868f
C1388 a_40868_n12168 a_40956_n12212 0.285629f
C1389 a_38292_n10980 VDD 0.244804f
C1390 a_44876_n14213 VDD 0.360805f
C1391 a_36140_n15348 a_36588_n15348 0.012001f
C1392 a_30676_n17252 VDD 0.212664f
C1393 a_47812_n20008 VDD 0.211703f
C1394 a_32909_841 a_31076_376 0.01529f
C1395 a_34895_376 a_35119_398 0.538085f
C1396 a_47924_n17252 a_47812_n18440 0.026657f
C1397 a_42324_n5896 a_41964_n5940 0.087174f
C1398 a_31324_n18484 a_31772_n18484 0.012882f
C1399 a_35268_n18440 a_35356_n18484 0.285629f
C1400 a_22052_n20008 a_21692_n20052 0.087066f
C1401 a_40196_n1884 VDD 0.460057f
C1402 a_25831_n11428 a_28335_n10644 0.010161f
C1403 a_38268_n9076 a_38380_n9509 0.026339f
C1404 a_41988_n20388 a_42436_n20388 0.013276f
C1405 a_41204_n4708 VDD 0.22954f
C1406 a_46108_n10644 a_46556_n10644 0.012552f
C1407 a_47812_n10600 a_47900_n10644 0.285629f
C1408 a_33832_n8572 VDD 0.47664f
C1409 a_46020_n12168 a_45660_n12212 0.086905f
C1410 a_41864_1394 a_42860_n101 0.0787f
C1411 a_32650_n12168 VDD 0.612661f
C1412 a_43108_n13736 a_43196_n13780 0.285629f
C1413 a_39164_n13780 a_39612_n13780 0.012882f
C1414 a_33252_n1192 a_33077_n1191 0.366162f
C1415 a_22052_n15304 VDD 0.204196f
C1416 a_43556_n15304 a_43196_n15348 0.087066f
C1417 a_22820_n2804 a_27672_n3543 0.012669f
C1418 a_22500_n1976 a_23319_n2759 0.022054f
C1419 a_25636_n18440 VDD 0.213265f
C1420 a_40956_n16916 a_41404_n16916 0.012882f
C1421 a_43868_n20485 VDD 0.362267f
C1422 a_38628_n18440 a_38268_n18484 0.087066f
C1423 a_46556_n5940 a_47004_n5940 0.012222f
C1424 a_28412_n20052 a_28860_n20052 0.012001f
C1425 a_45684_n4 a_45572_n1192 0.026657f
C1426 a_23507_n2759 VDD 0.609832f
C1427 a_47452_n9076 a_47564_n9509 0.026339f
C1428 a_31235_n9860 a_29992_n11150 0.229423f
C1429 a_29612_n8292 VDD 1.48038f
C1430 a_28927_n10160 a_31279_n11728 0.013151f
C1431 a_29332_n11301 a_30604_n11029 0.05539f
C1432 a_22220_n12996 a_21892_n12952 0.522083f
C1433 a_25724_n14564 a_25831_n12996 0.025245f
C1434 a_47364_n9032 VDD 0.205948f
C1435 a_25831_n12996 a_27639_n12537 0.024481f
C1436 a_41852_n12212 a_41740_n12645 0.026339f
C1437 a_38716_n12212 VDD 0.323196f
C1438 a_21772_n12996 a_23564_n20836 0.04672f
C1439 a_38628_n15304 VDD 0.214363f
C1440 a_47004_n15348 a_47452_n15348 0.012222f
C1441 a_32860_n2020 a_33120_n3884 0.017787f
C1442 a_33564_n18484 VDD 0.315469f
C1443 a_21692_2431 a_22052_1944 0.287426f
C1444 a_21604_n5067 a_22444_n5156 0.010538f
C1445 a_45124_376 a_45572_376 0.013276f
C1446 a_44452_n20388 VDD 0.23096f
C1447 a_45124_n18440 a_45572_n18440 0.013276f
C1448 a_34460_n18484 a_34348_n18917 0.026339f
C1449 a_29559_n6456 a_29123_n6679 0.01453f
C1450 a_35716_n20008 a_35356_n20052 0.087066f
C1451 a_23564_n8292 a_23816_n8544 0.038606f
C1452 a_47564_n7941 a_48012_n7941 0.012882f
C1453 a_42436_n2760 VDD 0.20462f
C1454 a_27516_n20052 XRST 0.025405f
C1455 a_28121_n10980 a_28300_n15348 0.062797f
C1456 a_25724_n14564 VDD 0.796932f
C1457 a_31760_n12168 a_31559_n13692 0.364366f
C1458 a_27639_n12537 VDD 0.803635f
C1459 a_22588_n15781 VDD 0.312053f
C1460 a_37452_n3888 a_37585_n3140 0.156824f
C1461 a_47364_n18440 VDD 0.205948f
C1462 a_21692_2431 a_26692_1564 0.016598f
C1463 a_38380_n17349 a_38828_n17349 0.012882f
C1464 a_28076_n17349 a_27988_n17252 0.285629f
C1465 a_45772_n6373 a_46220_n6373 0.012882f
C1466 a_40396_n6373 a_40308_n6276 0.285629f
C1467 a_41404_n18484 a_41292_n18917 0.026339f
C1468 a_42212_n20008 a_42660_n20008 0.013276f
C1469 a_38628_n20008 a_38716_n20052 0.285629f
C1470 a_37396_n9412 a_37844_n9412 0.013276f
C1471 a_45324_n9509 a_45236_n9412 0.285629f
C1472 a_25831_n11428 a_24684_n16432 0.51496f
C1473 a_40196_1944 VDD 0.867222f
C1474 a_48012_n6373 VDD 0.343411f
C1475 a_43980_n11077 a_43892_n10980 0.285629f
C1476 a_27281_n16854 a_27526_n13714 0.051134f
C1477 a_23564_n8292 a_24116_n15216 0.027664f
C1478 a_39636_n9412 VDD 0.209407f
C1479 a_37708_n12645 a_38068_n12548 0.086905f
C1480 a_25831_n12996 a_25237_n13735 0.054353f
C1481 a_46668_n12645 a_47116_n12645 0.012882f
C1482 a_33900_n14213 a_34260_n14116 0.087066f
C1483 a_29560_n3544 a_31248_n3544 0.012396f
C1484 a_37932_n15781 a_37844_n15684 0.285629f
C1485 a_46220_n15781 a_46668_n15781 0.012882f
C1486 a_24631_n3588 a_31392_n2760 0.51625f
C1487 a_26796_1515 a_27736_1248 0.056721f
C1488 a_25936_1564 a_28048_1248 0.277491f
C1489 a_39276_n18917 VDD 0.320362f
C1490 a_39612_n4805 a_40060_n4805 0.012222f
C1491 a_38828_n17349 a_39188_n17252 0.087066f
C1492 a_23484_n18917 a_23844_n18820 0.087174f
C1493 a_37036_n18917 a_37484_n18917 0.012882f
C1494 a_26531_n8639 a_26861_n8567 0.538085f
C1495 a_38068_n7844 a_38180_n9032 0.026657f
C1496 a_22568_n8944 a_22772_n8944 0.66083f
C1497 a_24233_n8684 a_21872_n9394 0.023272f
C1498 a_46668_n3237 VDD 0.318516f
C1499 a_29532_n10311 a_30599_n12167 0.017506f
C1500 a_21772_n9860 a_24964_n14116 0.844873f
C1501 a_32158_n12212 a_32650_n12168 0.086963f
C1502 a_46580_n10980 a_47028_n10980 0.013276f
C1503 a_31460_n10116 VDD 1.8252f
C1504 a_25237_n13735 VDD 0.502736f
C1505 a_36388_n1572 a_38312_n1975 0.013065f
C1506 a_36052_n14116 a_36500_n14116 0.013276f
C1507 a_44876_n14213 a_44788_n14116 0.285629f
C1508 a_22588_n16916 VDD 0.312663f
C1509 a_25237_n4327 a_28144_n4708 0.023385f
C1510 a_44428_n3237 a_44876_n3237 0.012882f
C1511 a_39948_n3237 a_39860_n3140 0.285629f
C1512 a_34471_1575 a_35064_1506 0.361958f
C1513 a_34260_n18820 VDD 0.206648f
C1514 a_44876_n4805 a_44788_n4708 0.285629f
C1515 a_39188_n17252 a_39636_n17252 0.013276f
C1516 a_25972_n6276 a_26643_n8292 0.01901f
C1517 a_34796_n18917 a_34708_n18820 0.285629f
C1518 a_30204_n20485 a_30652_n20485 0.013103f
C1519 a_28927_n10160 a_29444_n10116 0.029788f
C1520 a_28492_332 VDD 0.939787f
C1521 a_42748_n7508 VDD 0.315469f
C1522 a_40532_n10980 a_40420_n12168 0.026657f
C1523 a_40508_n10644 VDD 0.313885f
C1524 a_22016_n13665 a_23816_n13248 0.510371f
C1525 a_38180_n13736 VDD 0.24541f
C1526 a_34953_n1572 a_34248_n3310 0.148368f
C1527 a_44764_n1669 a_44676_n1572 0.285629f
C1528 a_39972_n16872 VDD 0.207295f
C1529 a_22052_n16872 a_22140_n16916 0.285629f
C1530 a_23396_n16872 a_23844_n16872 0.013276f
C1531 a_43416_1248 a_43728_1248 0.119687f
C1532 a_27428_n20008 VDD 0.206367f
C1533 a_33812_n17252 a_33924_n18440 0.026657f
C1534 a_24672_n11339 a_25524_n6635 0.021654f
C1535 a_45324_n18917 a_45684_n18820 0.087066f
C1536 a_31796_n18820 a_32244_n18820 0.013276f
C1537 a_33077_n1191 VDD 0.603685f
C1538 a_30652_n20485 a_30564_n20388 0.285629f
C1539 a_42212_n9032 a_42660_n9032 0.013276f
C1540 a_26531_n8639 a_26266_n9240 0.01478f
C1541 a_38628_n9032 a_38268_n9076 0.087066f
C1542 a_39308_n452 VDD 0.389039f
C1543 a_42748_n4372 VDD 0.315559f
C1544 a_38951_420 VDD 0.806241f
C1545 a_25020_n11383 a_30604_n11029 0.029899f
C1546 VDD CLK 3.7927f
C1547 a_38604_n7941 VDD 0.322493f
C1548 a_47028_n10980 a_46916_n12168 0.026657f
C1549 a_30092_n10980 VDD 0.010384f
C1550 a_43444_n12548 a_43556_n13736 0.026657f
C1551 a_41652_n14116 a_41764_n15304 0.026657f
C1552 a_29420_n17349 VDD 0.328085f
C1553 a_30788_n16872 a_30428_n16916 0.087174f
C1554 a_44340_n15684 a_44452_n16872 0.026657f
C1555 a_35849_n1192 a_35816_n174 0.427968f
C1556 a_33564_n20052 VDD 0.296789f
C1557 a_27628_n18484 a_28076_n18484 0.012552f
C1558 a_40508_n7508 a_40956_n7508 0.012882f
C1559 a_28660_n18820 a_28772_n20008 0.026657f
C1560 a_44452_n7464 a_44540_n7508 0.285629f
C1561 a_25647_n1976 VDD 0.764014f
C1562 a_30564_n20388 a_31012_n20388 0.013276f
C1563 a_25831_n11428 a_28624_n9394 0.396836f
C1564 a_41628_n20485 a_41988_n20388 0.087174f
C1565 a_38268_n10644 a_38716_n10644 0.012882f
C1566 a_42212_n10600 a_42300_n10644 0.285629f
C1567 a_28927_n10160 a_29744_n10980 0.014921f
C1568 a_29444_n10116 a_29332_n11301 0.030345f
C1569 a_46580_n7844 VDD 0.209016f
C1570 a_28009_n12168 a_27744_n12908 0.108149f
C1571 a_40868_n12168 a_40508_n12212 0.087066f
C1572 a_37844_n10980 VDD 0.215049f
C1573 a_35692_n13780 a_36140_n13780 0.012552f
C1574 a_34271_376 a_34068_n4 0.023823f
C1575 a_44428_n14213 VDD 0.321554f
C1576 a_30228_n17252 VDD 0.210675f
C1577 a_37732_n16872 a_38180_n16872 0.013276f
C1578 a_32579_769 a_31076_376 0.013404f
C1579 a_47364_n20008 VDD 0.205948f
C1580 a_35268_n18440 a_34908_n18484 0.087066f
C1581 a_23816_n5408 a_24573_n6724 0.022382f
C1582 a_41876_n5896 a_41964_n5940 0.285629f
C1583 a_22712_n7420 a_22876_n8988 0.019191f
C1584 a_35604_n18820 a_35716_n20008 0.026657f
C1585 a_21604_n20008 a_21692_n20052 0.285629f
C1586 a_38716_n7508 a_38604_n7941 0.026339f
C1587 a_25188_n20008 a_25636_n20008 0.013276f
C1588 a_37221_n3543 VDD 1.3222f
C1589 a_25642_n9816 a_26266_n9240 0.107109f
C1590 a_40420_n4708 VDD 0.211862f
C1591 a_47812_n10600 a_47452_n10644 0.086635f
C1592 a_46916_n12168 a_47364_n12168 0.013276f
C1593 a_45572_n12168 a_45660_n12212 0.285629f
C1594 a_32026_n12168 VDD 0.705154f
C1595 a_41864_1394 a_42412_n101 0.031841f
C1596 a_43108_n13736 a_42748_n13780 0.087066f
C1597 a_31656_n704 a_33077_n1191 0.016173f
C1598 a_21604_n15304 VDD 0.224005f
C1599 a_43108_n15304 a_43196_n15348 0.285629f
C1600 a_39164_n15348 a_39612_n15348 0.012882f
C1601 a_37785_n364 a_37680_n320 0.116059f
C1602 a_25188_n18440 VDD 0.217152f
C1603 a_38295_332 a_37368_n320 0.018241f
C1604 a_40508_n4372 a_40956_n4372 0.013103f
C1605 a_32668_n16916 a_32556_n17349 0.026339f
C1606 a_24631_n3588 a_24492_n5156 0.018971f
C1607 a_43420_n20485 VDD 0.332331f
C1608 a_41764_n18440 a_42212_n18440 0.013276f
C1609 a_38180_n18440 a_38268_n18484 0.285629f
C1610 a_42548_n18820 a_42660_n20008 0.026657f
C1611 a_47900_n7508 a_48012_n7941 0.026339f
C1612 a_36364_n7941 a_36812_n7941 0.013103f
C1613 a_30472_n9815 a_29992_n11150 0.096849f
C1614 a_25831_n11428 a_25500_n10644 0.013083f
C1615 a_35568_n4 VDD 0.810261f
C1616 a_29332_n11301 a_29744_n10980 0.536965f
C1617 a_46916_n9032 VDD 0.205962f
C1618 a_25831_n12996 a_25132_n16432 1.02164f
C1619 a_26239_n12996 a_25559_n12548 0.188134f
C1620 a_26563_n12212 a_27526_n13714 0.048456f
C1621 a_38268_n12212 VDD 0.358365f
C1622 a_46556_n13780 a_47004_n13780 0.012222f
C1623 a_38180_n15304 VDD 0.245127f
C1624 a_30555_n2729 a_29560_n3544 0.023304f
C1625 a_43420_n2804 a_43868_n2804 0.013103f
C1626 a_37372_n15348 a_37484_n15781 0.026339f
C1627 a_27988_n4328 a_28225_n4327 0.059868f
C1628 a_21692_2431 a_21604_2475 0.508857f
C1629 a_33116_n18484 VDD 0.332191f
C1630 a_39612_n16916 a_39724_n17349 0.026339f
C1631 a_43780_n20388 VDD 0.213385f
C1632 a_29559_n6456 a_30320_n6636 0.042802f
C1633 a_46108_n5940 a_46220_n6373 0.026339f
C1634 a_29211_n6724 a_29123_n6679 0.121284f
C1635 a_42548_n7844 CLK 0.029747f
C1636 a_35268_n20008 a_35356_n20052 0.285629f
C1637 a_31324_n20052 a_31772_n20052 0.012882f
C1638 a_40396_n7941 a_40308_n7844 0.285629f
C1639 a_41988_n2760 VDD 0.204447f
C1640 a_29992_n11150 a_28335_n10644 0.032527f
C1641 a_41740_n9509 a_42188_n9509 0.012882f
C1642 a_35468_n12645 a_35916_n12645 0.013103f
C1643 a_31760_n12168 a_31664_n13292 0.103816f
C1644 a_25132_n16432 VDD 0.629585f
C1645 a_22918_n2020 a_23542_n1754 0.106585f
C1646 a_21916_n1975 a_25647_n1976 0.031661f
C1647 a_31459_n14564 a_31789_n14564 0.538085f
C1648 a_22140_n15781 VDD 0.296789f
C1649 a_37452_n3888 a_22052_n4708 0.059876f
C1650 a_35244_n15781 a_35692_n15781 0.012882f
C1651 a_23507_n2759 a_26047_n4328 0.054584f
C1652 a_46556_n15348 a_46668_n15781 0.026339f
C1653 a_25759_n3544 a_26383_n2968 0.104193f
C1654 a_28736_1944 a_25600_n5895 0.052833f
C1655 a_21692_2431 a_26488_1564 0.027059f
C1656 a_46916_n18440 VDD 0.205962f
C1657 a_26060_n18917 a_26508_n18917 0.012882f
C1658 a_39948_n6373 a_40308_n6276 0.086635f
C1659 a_38628_n20008 a_38268_n20052 0.087066f
C1660 a_44340_n7844 a_44788_n7844 0.013276f
C1661 a_27932_n3543 VDD 0.319149f
C1662 a_44876_n9509 a_45236_n9412 0.087066f
C1663 a_25831_n11428 a_25559_n10980 0.058436f
C1664 a_47564_n6373 VDD 0.315469f
C1665 a_43532_n11077 a_43892_n10980 0.087066f
C1666 a_27281_n16854 a_27302_n13160 0.044784f
C1667 a_39188_n9412 VDD 0.211136f
C1668 a_23564_n11428 a_25160_n14816 0.034774f
C1669 a_37708_n12645 a_37620_n12548 0.285629f
C1670 a_46580_n4 a_46468_n1192 0.026657f
C1671 a_33900_n14213 a_33812_n14116 0.285629f
C1672 a_42188_n14213 a_42636_n14213 0.012882f
C1673 a_48012_n15781 VDD 0.343411f
C1674 a_34000_n3140 a_36112_n3456 0.277491f
C1675 a_37484_n15781 a_37844_n15684 0.087066f
C1676 a_29560_n3544 a_30820_n3544 0.012072f
C1677 a_34552_n3140 a_34756_n3140 0.66083f
C1678 a_47900_n2804 a_48012_n3237 0.026339f
C1679 a_42604_n2020 a_46580_n4 0.012286f
C1680 a_24631_n3588 a_31412_n2276 0.525637f
C1681 a_42604_n2020 a_46108_n1669 0.017891f
C1682 a_26284_1564 a_26488_1564 0.048436f
C1683 a_26796_1515 a_26692_1564 0.026665f
C1684 a_38828_n18917 VDD 0.322604f
C1685 a_25936_1564 a_28153_1204 0.020455f
C1686 a_27988_n17252 a_28436_n17252 0.013276f
C1687 a_38828_n17349 a_38740_n17252 0.285629f
C1688 a_23484_n18917 a_23396_n18820 0.285629f
C1689 a_45684_n6276 a_46132_n6276 0.013276f
C1690 a_42748_n9076 CLK 0.012909f
C1691 a_36252_n20052 a_36252_n20485 0.05841f
C1692 a_45124_n20008 a_45572_n20008 0.013276f
C1693 a_23564_n8292 a_24965_n9860 1.82382f
C1694 a_42660_n12168 CLK 0.017841f
C1695 a_46220_n3237 VDD 0.320246f
C1696 a_28335_n10644 a_28247_n10599 0.081541f
C1697 a_22264_n8988 a_22700_n12080 0.019845f
C1698 a_35324_1564 VDD 0.298894f
C1699 a_32158_n12212 a_32026_n12168 0.484914f
C1700 a_30136_n10600 VDD 0.259016f
C1701 a_39412_n12548 a_39860_n12548 0.013276f
C1702 a_23816_n13248 VDD 1.38103f
C1703 a_44428_n14213 a_44788_n14116 0.087066f
C1704 a_36388_n1572 a_37632_n2020 0.55986f
C1705 a_22500_n1976 a_22016_n1121 0.048337f
C1706 a_22140_n16916 VDD 0.312663f
C1707 a_39500_n3237 a_39860_n3140 0.086742f
C1708 a_39636_n15684 a_40084_n15684 0.013276f
C1709 a_22500_n1976 a_23004_n2332 1.75958f
C1710 a_33812_n18820 VDD 0.206648f
C1711 a_34576_1204 a_34872_1619 0.05539f
C1712 a_44428_n4805 a_44788_n4708 0.087066f
C1713 a_38180_n4708 a_38628_n4708 0.013276f
C1714 a_41652_n6276 a_41764_n7464 0.026657f
C1715 a_34348_n18917 a_34708_n18820 0.087066f
C1716 a_47564_n18917 a_48012_n18917 0.012882f
C1717 a_27540_n3797 VDD 0.475465f
C1718 a_41652_n9412 a_41764_n10600 0.026657f
C1719 a_27572_860 VDD 0.482724f
C1720 a_42300_n7508 VDD 0.315469f
C1721 a_42748_n18484 CLK 0.012909f
C1722 a_40060_n10644 VDD 0.314419f
C1723 a_21604_n13252 a_23816_n13248 0.042802f
C1724 a_22016_n13665 a_24233_n13388 0.020455f
C1725 a_37732_n13736 VDD 0.213395f
C1726 a_44316_n1669 a_44676_n1572 0.087174f
C1727 a_46580_n14116 a_47028_n14116 0.013276f
C1728 a_33812_n14116 a_33812_n15304 0.05841f
C1729 a_39524_n16872 VDD 0.209499f
C1730 a_22052_n16872 a_21692_n16916 0.086905f
C1731 a_46132_n3140 a_46580_n3140 0.013276f
C1732 a_26980_n20008 VDD 0.206367f
C1733 a_43416_1248 a_43833_1204 0.633318f
C1734 a_37859_377 a_30104_n1148 0.017428f
C1735 a_22948_n18440 a_23396_n18440 0.013276f
C1736 a_24672_n11339 a_25612_n6679 0.013902f
C1737 a_37284_n7464 a_37732_n7464 0.013276f
C1738 a_45324_n18917 a_45236_n18820 0.285629f
C1739 a_30612_n1104 VDD 0.299323f
C1740 a_38180_n9032 a_38268_n9076 0.285629f
C1741 a_41180_n20485 a_41628_n20485 0.013103f
C1742 a_30204_n20485 a_30564_n20388 0.087174f
C1743 a_42300_n4372 VDD 0.315559f
C1744 a_25020_n11383 a_29744_n10980 0.044096f
C1745 a_39056_820 VDD 1.80728f
C1746 a_38156_n7941 VDD 0.355226f
C1747 a_30604_n11029 VDD 0.261506f
C1748 a_32412_n13648 VDD 0.301311f
C1749 a_21716_n2229 a_22164_n2760 0.195633f
C1750 a_28972_n17349 VDD 0.327647f
C1751 a_27988_n20388 a_27988_n18440 0.018105f
C1752 a_33476_n16872 a_33924_n16872 0.013276f
C1753 a_42100_n3140 a_42212_n4328 0.026657f
C1754 a_30340_n16872 a_30428_n16916 0.285629f
C1755 a_33116_n20052 VDD 0.298821f
C1756 a_40532_n17252 a_40420_n18440 0.026657f
C1757 a_42548_n18820 a_42996_n18820 0.013276f
C1758 a_44452_n7464 a_44092_n7508 0.086635f
C1759 a_25972_n6276 a_21872_n9394 0.015084f
C1760 a_24315_n2759 VDD 0.68751f
C1761 a_41628_n20485 a_41540_n20388 0.285629f
C1762 a_25831_n11428 a_29800_n9815 0.014829f
C1763 a_44540_n9076 a_45124_n9032 0.016748f
C1764 a_27414_n5112 VDD 0.327345f
C1765 a_42212_n10600 a_41852_n10644 0.087066f
C1766 a_42948_n1976 a_42884_n1192 0.050489f
C1767 a_46132_n7844 VDD 0.210512f
C1768 a_24684_n16432 a_25642_n13736 0.011212f
C1769 a_40420_n12168 a_40508_n12212 0.285629f
C1770 a_37396_n10980 VDD 0.212402f
C1771 a_40260_n408 a_42948_n1976 0.059024f
C1772 a_27055_n1192 a_27279_n1170 0.538085f
C1773 a_34403_332 a_34068_n4 0.223963f
C1774 a_43980_n14213 VDD 0.31896f
C1775 a_35692_n15348 a_36140_n15348 0.013103f
C1776 a_29780_n17252 VDD 0.209282f
C1777 a_22052_n4708 a_28548_n5112 0.012902f
C1778 a_34271_376 a_34895_376 0.104193f
C1779 a_46916_n20008 VDD 0.205962f
C1780 a_30876_n18484 a_31324_n18484 0.012882f
C1781 a_41876_n5896 a_41516_n5940 0.087174f
C1782 a_34820_n18440 a_34908_n18484 0.285629f
C1783 a_47476_n17252 a_47364_n18440 0.026657f
C1784 a_33497_n9032 a_29532_n10311 0.035196f
C1785 a_22712_n7420 a_22264_n8988 0.02881f
C1786 a_39648_n2020 VDD 0.456298f
C1787 a_37820_n9076 a_37932_n9509 0.026339f
C1788 a_41540_n20388 a_41988_n20388 0.013276f
C1789 a_25237_n10599 a_26266_n9240 0.055668f
C1790 a_39972_n4708 VDD 0.207445f
C1791 a_45660_n10644 a_46108_n10644 0.012552f
C1792 a_47364_n10600 a_47452_n10644 0.285629f
C1793 a_45572_n12168 a_45212_n12212 0.086905f
C1794 a_31279_n11728 VDD 0.637768f
C1795 a_32073_n844 a_33077_n1191 0.111715f
C1796 a_30159_n13296 a_31789_n14564 0.016087f
C1797 a_38716_n13780 a_39164_n13780 0.012882f
C1798 a_42660_n13736 a_42748_n13780 0.285629f
C1799 a_34248_n3310 a_34348_n3140 0.092119f
C1800 a_43108_n15304 a_42748_n15348 0.087066f
C1801 a_27988_n20388 a_26755_n16132 0.045856f
C1802 a_38733_n2295 a_39357_n2228 0.104193f
C1803 a_32984_n2672 a_33188_n2672 0.66083f
C1804 a_22820_n2804 a_26383_n2968 0.013488f
C1805 a_37368_n320 a_37680_n320 0.119687f
C1806 a_24740_n18440 VDD 0.242651f
C1807 a_44452_n16872 a_44540_n16916 0.285629f
C1808 a_40508_n16916 a_40956_n16916 0.012882f
C1809 a_44452_n4328 a_44540_n4372 0.285629f
C1810 a_42972_n20485 VDD 0.329322f
C1811 a_38180_n18440 a_37820_n18484 0.087066f
C1812 a_47812_n5896 a_47900_n5940 0.285629f
C1813 a_46108_n5940 a_46556_n5940 0.012552f
C1814 a_27964_n20052 a_28412_n20052 0.012882f
C1815 a_24403_n2414 VDD 0.726292f
C1816 a_30472_n9815 a_25724_n14564 0.194615f
C1817 a_35156_n325 a_35119_n1170 0.035793f
C1818 a_47004_n9076 a_47116_n9509 0.026339f
C1819 a_35156_n325 a_37785_n364 0.019043f
C1820 a_25412_n5895 VDD 0.596387f
C1821 a_28927_n10160 a_29540_n11728 0.036041f
C1822 a_46468_n9032 VDD 0.209055f
C1823 a_41404_n12212 a_41292_n12645 0.026339f
C1824 a_26983_n12728 a_27744_n12908 0.042802f
C1825 a_26563_n12212 a_27302_n13160 0.064633f
C1826 a_25831_n12996 a_25559_n12548 0.02258f
C1827 a_37820_n12212 VDD 0.324562f
C1828 a_37732_n15304 VDD 0.213126f
C1829 a_32860_n2020 a_32359_n4372 0.022396f
C1830 a_46556_n15348 a_47004_n15348 0.012222f
C1831 a_32668_n18484 VDD 0.317969f
C1832 a_43332_n20388 VDD 0.205276f
C1833 a_44540_332 a_45124_376 0.016748f
C1834 a_44540_n18484 a_45124_n18440 0.016748f
C1835 a_29211_n6724 a_30320_n6636 0.019043f
C1836 a_34012_n18484 a_33900_n18917 0.026339f
C1837 a_25612_n6679 a_30740_n7464 0.030106f
C1838 a_42100_n7844 CLK 0.023004f
C1839 a_35268_n20008 a_34908_n20052 0.087066f
C1840 a_47116_n7941 a_47564_n7941 0.012882f
C1841 a_39948_n7941 a_40308_n7844 0.086742f
C1842 a_41540_n2760 VDD 0.207105f
C1843 a_24965_n9860 a_22016_n10529 0.044092f
C1844 a_47900_n5940 VDD 0.335152f
C1845 a_30871_n11728 a_35804_n12212 0.025595f
C1846 a_40172_n11077 a_40620_n11077 0.012222f
C1847 a_25559_n12548 VDD 0.963766f
C1848 a_42748_n20052 CLK 0.012909f
C1849 a_31459_n14564 a_28752_n15348 0.03379f
C1850 a_21916_n1975 a_24315_n2759 0.036608f
C1851 a_21692_n15781 VDD 0.300735f
C1852 a_23507_n2759 a_25423_n4328 0.465142f
C1853 a_25237_n4327 a_26383_n2968 0.064141f
C1854 a_26607_1966 a_25524_1243 0.031731f
C1855 a_46468_n18440 VDD 0.209055f
C1856 a_24604_n17349 a_24516_n17252 0.285629f
C1857 a_37932_n17349 a_38380_n17349 0.012882f
C1858 a_39948_n6373 a_39860_n6276 0.285629f
C1859 a_45324_n6373 a_45772_n6373 0.012882f
C1860 a_38180_n20008 a_38268_n20052 0.285629f
C1861 a_41764_n20008 a_42212_n20008 0.013276f
C1862 a_27672_n3543 VDD 0.459055f
C1863 a_36948_n9412 a_37396_n9412 0.013276f
C1864 a_44876_n9509 a_44788_n9412 0.285629f
C1865 a_47476_n4 a_47924_n4 0.013276f
C1866 a_47116_n6373 VDD 0.315469f
C1867 a_43532_n11077 a_43444_n10980 0.285629f
C1868 a_38740_n9412 VDD 0.213797f
C1869 a_37260_n12645 a_37620_n12548 0.086905f
C1870 a_46220_n12645 a_46668_n12645 0.012882f
C1871 a_48012_n12645 VDD 0.343411f
C1872 a_33452_n14213 a_33812_n14116 0.087066f
C1873 a_47564_n15781 VDD 0.315469f
C1874 a_45772_n15781 a_46220_n15781 0.012882f
C1875 a_37484_n15781 a_37396_n15684 0.285629f
C1876 a_34860_n3189 a_35800_n3456 0.056721f
C1877 a_29560_n3544 a_30616_n3544 0.011094f
C1878 a_34000_n3140 a_36217_n3500 0.020455f
C1879 a_24631_n3588 a_30555_n2729 0.029185f
C1880 a_42604_n2020 a_45660_n1669 0.017213f
C1881 a_25936_1564 a_27736_1248 0.510371f
C1882 a_26796_1515 a_26488_1564 0.934191f
C1883 a_38380_n18917 VDD 0.342527f
C1884 a_35816_n174 a_35568_n4 0.355778f
C1885 a_39164_n4805 a_39612_n4805 0.012552f
C1886 a_38380_n17349 a_38740_n17252 0.087066f
C1887 a_36588_n18917 a_37036_n18917 0.012882f
C1888 a_23036_n18917 a_23396_n18820 0.087174f
C1889 a_42300_n9076 CLK 0.048577f
C1890 a_22876_n8988 a_22772_n8944 0.026665f
C1891 a_37620_n7844 a_37732_n9032 0.026657f
C1892 a_45772_n3237 VDD 0.322355f
C1893 a_42212_n12168 CLK 0.037136f
C1894 a_28335_n10644 a_31460_n10116 0.02173f
C1895 a_34872_1619 VDD 0.244331f
C1896 a_27540_n20747 XRST 0.743784f
C1897 a_30036_n7464 VDD 0.605932f
C1898 a_46132_n10980 a_46580_n10980 0.013276f
C1899 a_29444_n10116 VDD 0.543173f
C1900 a_24233_n13388 VDD 0.508785f
C1901 a_44428_n14213 a_44340_n14116 0.285629f
C1902 a_35604_n14116 a_36052_n14116 0.013276f
C1903 a_22500_n1976 a_21604_n708 0.017215f
C1904 a_21692_n16916 VDD 0.317437f
C1905 a_39500_n3237 a_39412_n3140 0.285629f
C1906 a_43980_n3237 a_44428_n3237 0.012882f
C1907 a_33815_1384 a_34872_1619 0.056721f
C1908 a_33364_n18820 VDD 0.227401f
C1909 a_38740_n17252 a_39188_n17252 0.013276f
C1910 a_44428_n4805 a_44340_n4708 0.285629f
C1911 a_34348_n18917 a_34260_n18820 0.285629f
C1912 a_28617_n8548 a_25831_n11428 0.986564f
C1913 a_29756_n20485 a_30204_n20485 0.013103f
C1914 a_28144_n4708 VDD 1.27369f
C1915 a_28927_n10160 a_28435_n10599 0.720338f
C1916 a_25724_n14564 a_24684_n16432 0.010715f
C1917 a_41852_n7508 VDD 0.315469f
C1918 a_40084_n10980 a_39972_n12168 0.026657f
C1919 a_39612_n10644 VDD 0.317476f
C1920 a_42300_n18484 CLK 0.048577f
C1921 a_22364_n13648 a_22568_n13648 0.048436f
C1922 a_21604_n13252 a_24233_n13388 0.019043f
C1923 a_37284_n13736 VDD 0.232558f
C1924 a_44316_n1669 a_44228_n1572 0.285629f
C1925 a_39076_n16872 VDD 0.211414f
C1926 a_36500_n15684 a_36612_n16872 0.026657f
C1927 a_21604_n16872 a_21692_n16916 0.285629f
C1928 a_22948_n16872 a_23396_n16872 0.013276f
C1929 a_26532_n20008 VDD 0.206917f
C1930 a_23228_n6679 a_23619_n6724 0.010772f
C1931 a_24672_n11339 a_24573_n6724 0.090347f
C1932 a_33364_n17252 a_33476_n18440 0.026657f
C1933 a_31348_n18820 a_31796_n18820 0.013276f
C1934 a_44876_n18917 a_45236_n18820 0.087066f
C1935 a_47476_n4 a_47364_n1192 0.026657f
C1936 a_31968_n704 VDD 0.025368f
C1937 a_38180_n9032 a_37820_n9076 0.087066f
C1938 a_41764_n9032 a_42212_n9032 0.013276f
C1939 a_30204_n20485 a_30116_n20388 0.285629f
C1940 a_41852_n4372 VDD 0.315559f
C1941 a_25020_n11383 a_28121_n10980 0.048028f
C1942 a_37708_n7941 VDD 0.322183f
C1943 a_46580_n10980 a_46468_n12168 0.026657f
C1944 a_29744_n10980 VDD 0.822366f
C1945 a_42996_n12548 a_43108_n13736 0.026657f
C1946 a_47900_n13780 VDD 0.335152f
C1947 a_41204_n14116 a_41316_n15304 0.026657f
C1948 a_22820_n2804 a_22164_n2760 0.206411f
C1949 a_28524_n17349 VDD 0.31407f
C1950 a_27988_n20388 a_27540_n18440 0.041636f
C1951 a_27988_n4328 a_25972_n6276 0.043774f
C1952 a_25600_n5895 a_26154_n4536 0.012701f
C1953 a_43892_n15684 a_44004_n16872 0.026657f
C1954 a_32668_n20052 VDD 0.333905f
C1955 a_27180_n18484 a_27628_n18484 0.012552f
C1956 a_44004_n7464 a_44092_n7508 0.285629f
C1957 a_28212_n18820 a_28324_n20008 0.026657f
C1958 a_30396_n7508 a_31341_n8292 0.013814f
C1959 a_40060_n7508 a_40508_n7508 0.012882f
C1960 a_24578_n2020 VDD 0.837992f
C1961 a_41180_n20485 a_41540_n20388 0.087174f
C1962 a_30116_n20388 a_30564_n20388 0.013276f
C1963 a_25831_n11428 a_27281_n16854 0.011988f
C1964 a_40652_n1572 a_45684_n4 0.029747f
C1965 a_27190_n5112 VDD 0.596541f
C1966 a_37820_n10644 a_38268_n10644 0.012882f
C1967 a_41764_n10600 a_41852_n10644 0.285629f
C1968 a_25020_n11383 a_33364_n11384 0.018526f
C1969 a_28437_n13705 a_28121_n10980 0.027806f
C1970 a_32262_n452 a_33508_n408 0.010837f
C1971 a_42948_n1976 a_42157_n660 0.020396f
C1972 a_45684_n7844 VDD 0.212747f
C1973 a_40420_n12168 a_40060_n12212 0.087066f
C1974 a_36948_n10980 VDD 0.213596f
C1975 a_23816_n704 a_24128_n704 0.119687f
C1976 a_35244_n13780 a_35692_n13780 0.012552f
C1977 a_43532_n14213 VDD 0.317216f
C1978 a_29332_n17252 VDD 0.206765f
C1979 a_37284_n16872 a_37732_n16872 0.013276f
C1980 a_46468_n20008 VDD 0.209055f
C1981 a_24631_n3588 a_31076_376 0.133903f
C1982 a_43644_n705 a_44452_376 0.024871f
C1983 a_34403_332 a_34895_376 0.081624f
C1984 a_41428_n5896 a_41516_n5940 0.285629f
C1985 a_34820_n18440 a_34460_n18484 0.087066f
C1986 a_37372_n5940 a_37820_n5940 0.012222f
C1987 a_24740_n20008 a_25188_n20008 0.013276f
C1988 a_38268_n7508 a_38156_n7941 0.026339f
C1989 a_22712_n7420 a_22016_n8961 0.028885f
C1990 a_35156_n18820 a_35268_n20008 0.026657f
C1991 a_38984_n1975 VDD 0.451402f
C1992 a_25237_n10599 a_25642_n9816 0.488306f
C1993 a_22116_n9412 a_21892_n9816 0.013419f
C1994 a_39524_n4708 VDD 0.209769f
C1995 a_47364_n10600 a_47004_n10644 0.086742f
C1996 a_28225_n9031 VDD 0.967739f
C1997 a_45124_n12168 a_45212_n12212 0.285629f
C1998 a_46468_n12168 a_46916_n12168 0.013276f
C1999 a_30159_n13296 a_28752_n15348 0.074593f
C2000 a_34895_n1192 a_35119_n1170 0.538085f
C2001 a_31656_n704 a_31968_n704 0.119687f
C2002 a_42660_n13736 a_42300_n13780 0.087066f
C2003 a_47924_n14116 VDD 0.21239f
C2004 a_42660_n15304 a_42748_n15348 0.285629f
C2005 a_22164_n2760 a_25237_n4327 1.71197f
C2006 a_38716_n15348 a_39164_n15348 0.012882f
C2007 a_37368_n320 a_37785_n364 0.633318f
C2008 a_24292_n18440 VDD 0.218083f
C2009 a_40060_n4372 a_40508_n4372 0.013103f
C2010 a_44452_n4328 a_44092_n4372 0.086635f
C2011 a_44452_n16872 a_44092_n16916 0.086635f
C2012 a_32220_n16916 a_32108_n17349 0.026339f
C2013 a_42524_n20485 VDD 0.329322f
C2014 a_41316_n18440 a_41764_n18440 0.013276f
C2015 a_37732_n18440 a_37820_n18484 0.285629f
C2016 a_47812_n5896 a_47452_n5940 0.086635f
C2017 a_47452_n7508 a_47564_n7941 0.026339f
C2018 a_42100_n18820 a_42212_n20008 0.026657f
C2019 a_35156_n325 a_34895_n1192 0.021138f
C2020 a_28624_n9394 a_25724_n14564 0.011465f
C2021 a_37844_1564 OUT[2] 0.012283f
C2022 a_35156_n325 a_37368_n320 0.042802f
C2023 a_25724_n14564 a_24573_n12996 0.019816f
C2024 a_27281_n16854 a_27535_n12493 0.015371f
C2025 a_44540_n10644 a_44428_n11077 0.026339f
C2026 a_27391_n11384 a_28121_n10980 0.240599f
C2027 a_46020_n9032 VDD 0.210736f
C2028 a_26635_n12996 a_27744_n12908 0.019043f
C2029 a_37372_n12212 VDD 0.326159f
C2030 a_21772_n12996 a_22052_n15684 0.049548f
C2031 a_47812_n13736 a_47900_n13780 0.285629f
C2032 a_46108_n13780 a_46556_n13780 0.012552f
C2033 a_37284_n15304 VDD 0.232289f
C2034 a_32860_n2020 a_31787_n3969 0.01575f
C2035 a_42972_n2804 a_43420_n2804 0.013103f
C2036 a_27988_n20388 a_23564_n17700 0.09415f
C2037 a_32220_n18484 VDD 0.320004f
C2038 a_39164_n16916 a_39276_n17349 0.026339f
C2039 a_42884_n20388 VDD 0.203482f
C2040 a_29211_n6724 a_29559_n6456 0.633318f
C2041 a_45660_n5940 a_45772_n6373 0.026339f
C2042 a_25972_n6276 a_29123_n6679 0.338512f
C2043 a_30876_n20052 a_31324_n20052 0.012882f
C2044 a_39948_n7941 a_39860_n7844 0.285629f
C2045 a_34820_n20008 a_34908_n20052 0.285629f
C2046 a_41092_n2760 VDD 0.206217f
C2047 a_41292_n9509 a_41740_n9509 0.012882f
C2048 a_24965_n9860 a_21604_n10116 0.010875f
C2049 a_22264_n10556 a_22364_n10512 0.084652f
C2050 a_47452_n5940 VDD 0.313885f
C2051 a_30871_n11728 a_35356_n12212 0.01798f
C2052 a_35020_n12645 a_35468_n12645 0.013103f
C2053 a_42300_n20052 CLK 0.048949f
C2054 a_27820_n16432 a_27852_n14990 0.358902f
C2055 a_21916_n1975 a_24578_n2020 0.03493f
C2056 a_47900_n15348 VDD 0.335152f
C2057 a_46108_n15348 a_46220_n15781 0.026339f
C2058 a_22164_n2760 a_24128_n3840 0.012204f
C2059 a_34796_n15781 a_35244_n15781 0.012882f
C2060 a_26383_1944 a_25524_1243 0.041412f
C2061 a_46020_n18440 VDD 0.210736f
C2062 a_21692_2431 a_26796_1515 0.018157f
C2063 a_40508_n18484 a_40620_n18917 0.026339f
C2064 a_25612_n18917 a_26060_n18917 0.012882f
C2065 a_39500_n6373 a_39860_n6276 0.086742f
C2066 a_38180_n20008 a_37820_n20052 0.087066f
C2067 a_43892_n7844 a_44340_n7844 0.013276f
C2068 a_26607_n3544 VDD 0.307525f
C2069 a_44428_n9509 a_44788_n9412 0.087066f
C2070 a_39748_2475 VDD 0.499331f
C2071 a_46668_n6373 VDD 0.318039f
C2072 a_33572_n10980 a_33364_n11384 0.013419f
C2073 a_43084_n11077 a_43444_n10980 0.087066f
C2074 a_38292_n9412 VDD 0.243753f
C2075 a_37260_n12645 a_37172_n12548 0.285629f
C2076 a_47564_n12645 VDD 0.315469f
C2077 a_33452_n14213 a_33364_n14116 0.285629f
C2078 a_41740_n14213 a_42188_n14213 0.012882f
C2079 a_47116_n15781 VDD 0.315469f
C2080 a_34000_n3140 a_35800_n3456 0.510371f
C2081 a_34860_n3189 a_34756_n3140 0.026665f
C2082 a_37036_n15781 a_37396_n15684 0.087066f
C2083 a_34348_n3140 a_34552_n3140 0.048436f
C2084 a_36120_n4 VDD 0.362528f
C2085 a_47452_n2804 a_47564_n3237 0.026339f
C2086 a_25600_n5895 a_22052_n4708 0.015858f
C2087 a_42604_n2020 a_45212_n1669 0.012889f
C2088 a_37932_n18917 VDD 0.327654f
C2089 a_38380_n17349 a_38292_n17252 0.285629f
C2090 a_23564_n20836 a_24292_n18820 0.017973f
C2091 a_45236_n6276 a_45684_n6276 0.013276f
C2092 a_23036_n18917 a_22948_n18820 0.285629f
C2093 a_41852_n9076 CLK 0.013107f
C2094 a_23564_n8292 a_23949_n9860 0.039281f
C2095 a_22568_n8944 a_21872_n9394 0.018252f
C2096 a_35804_n20052 a_35804_n20485 0.05841f
C2097 a_44540_n20052 a_45124_n20008 0.016748f
C2098 a_45324_n3237 VDD 0.325321f
C2099 a_28335_n10644 a_30136_n10600 0.020642f
C2100 a_25020_n11383 a_28435_n10599 0.078502f
C2101 a_21772_n9860 a_23564_n11428 0.01446f
C2102 a_23479_n5156 a_25577_n14956 0.013277f
C2103 a_22264_n8988 a_22600_n12124 1.39342f
C2104 a_47476_n9412 a_47924_n9412 0.013276f
C2105 a_34367_1619 VDD 0.022335f
C2106 a_26844_n20485 XRST 0.048835f
C2107 a_30396_n7508 VDD 0.654923f
C2108 a_38964_n12548 a_39412_n12548 0.013276f
C2109 a_36744_n1954 a_36388_n1572 0.579288f
C2110 a_43980_n14213 a_44340_n14116 0.087066f
C2111 a_28548_n16872 VDD 0.133407f
C2112 a_39188_n15684 a_39636_n15684 0.013276f
C2113 a_48012_n15781 a_47924_n15684 0.285629f
C2114 a_33815_1384 a_34367_1619 0.119687f
C2115 a_34576_1204 a_35064_1506 0.08126f
C2116 a_32692_n18820 VDD 0.216918f
C2117 a_43980_n4805 a_44340_n4708 0.087066f
C2118 a_33900_n18917 a_34260_n18820 0.087066f
C2119 a_41204_n6276 a_41316_n7464 0.026657f
C2120 a_47116_n18917 a_47564_n18917 0.012882f
C2121 a_27988_n4328 a_30599_n12167 0.07614f
C2122 a_41204_n9412 a_41316_n10600 0.026657f
C2123 a_28437_n13705 a_28435_n10599 0.540581f
C2124 a_26756_n20388 XRST 0.013113f
C2125 a_41404_n7508 VDD 0.315469f
C2126 a_24684_n16432 a_25132_n16432 0.152985f
C2127 a_39164_n10644 VDD 0.319301f
C2128 a_41852_n18484 CLK 0.013107f
C2129 a_22876_n13692 a_22568_n13648 0.934191f
C2130 a_36588_n13780 VDD 0.321045f
C2131 a_33364_n14116 a_33364_n15304 0.05841f
C2132 a_46132_n14116 a_46580_n14116 0.013276f
C2133 a_43868_n1669 a_44228_n1572 0.087174f
C2134 a_38628_n16872 VDD 0.214363f
C2135 a_45684_n3140 a_46132_n3140 0.013276f
C2136 a_26084_n20008 VDD 0.209243f
C2137 a_23228_n6679 a_22968_n6679 0.509297f
C2138 a_24492_n5156 a_25612_n6679 0.219546f
C2139 a_22500_n18440 a_22948_n18440 0.013276f
C2140 a_22444_n5156 a_25972_n6276 0.048401f
C2141 a_44876_n18917 a_44788_n18820 0.285629f
C2142 a_40732_n20485 a_41180_n20485 0.013103f
C2143 a_37732_n9032 a_37820_n9076 0.285629f
C2144 a_21872_n9394 a_22264_n10556 0.040203f
C2145 a_29756_n20485 a_30116_n20388 0.087174f
C2146 a_41404_n4372 VDD 0.315559f
C2147 a_30871_n11728 a_33900_n11428 0.522567f
C2148 a_21772_n9860 a_22600_n12124 0.02796f
C2149 a_38295_332 VDD 1.35484f
C2150 a_37260_n7941 VDD 0.319373f
C2151 a_28121_n10980 VDD 0.832855f
C2152 a_47452_n13780 VDD 0.313885f
C2153 a_21692_2431 a_29295_n1400 0.055047f
C2154 a_28076_n17349 VDD 0.332877f
C2155 a_41652_n3140 a_41764_n4328 0.026657f
C2156 a_25600_n5895 a_25530_n5112 0.073571f
C2157 a_33028_n16872 a_33476_n16872 0.013276f
C2158 a_24913_864 a_25817_804 0.514036f
C2159 a_32220_n20052 VDD 0.335021f
C2160 a_40084_n17252 a_39972_n18440 0.026657f
C2161 a_30396_n7508 a_30676_n7844 0.148917f
C2162 a_44004_n7464 a_43644_n7508 0.087066f
C2163 a_42100_n18820 a_42548_n18820 0.013276f
C2164 a_23954_n2020 VDD 0.609394f
C2165 a_41180_n20485 a_41092_n20388 0.285629f
C2166 a_44092_n9076 a_44540_n9076 0.012001f
C2167 a_41764_n10600 a_41404_n10644 0.087066f
C2168 a_45236_n7844 VDD 0.229781f
C2169 a_26563_n12212 a_27535_n12493 0.049361f
C2170 a_44004_n12168 a_44452_n12168 0.013276f
C2171 a_39972_n12168 a_40060_n12212 0.285629f
C2172 a_33364_n11384 VDD 0.855405f
C2173 a_21772_n12996 a_23608_n15260 0.010392f
C2174 a_24233_n844 a_24128_n704 0.116059f
C2175 a_26431_n1192 a_27055_n1192 0.104193f
C2176 a_21692_2431 a_26631_7 0.017162f
C2177 a_43084_n14213 VDD 0.313885f
C2178 a_47924_n14116 a_47812_n15304 0.026657f
C2179 a_35244_n15348 a_35692_n15348 0.013103f
C2180 a_28884_n17252 VDD 0.209253f
C2181 a_30372_376 a_31076_376 0.223141f
C2182 a_46020_n20008 VDD 0.210736f
C2183 a_34403_332 a_34271_376 0.48859f
C2184 a_43644_n705 a_40260_n408 0.037233f
C2185 a_34372_n18440 a_34460_n18484 0.285629f
C2186 a_47028_n17252 a_46916_n18440 0.026657f
C2187 a_41428_n5896 a_41068_n5940 0.087174f
C2188 a_30428_n18484 a_30876_n18484 0.012882f
C2189 a_22712_n7420 a_21604_n8548 0.015849f
C2190 a_47452_n7508 a_47900_n7508 0.012001f
C2191 a_38312_n1975 VDD 0.490948f
C2192 a_42660_n10600 CLK 0.017841f
C2193 a_41092_n20388 a_41540_n20388 0.013276f
C2194 a_37372_n9076 a_37484_n9509 0.026339f
C2195 a_39076_n4708 VDD 0.214403f
C2196 a_45212_n10644 a_45660_n10644 0.012552f
C2197 a_46916_n10600 a_47004_n10644 0.285629f
C2198 a_28927_n10160 a_28300_n15348 0.212614f
C2199 a_29540_n11728 VDD 0.567455f
C2200 a_42212_n13736 a_42300_n13780 0.285629f
C2201 a_32073_n844 a_31968_n704 0.116059f
C2202 a_38268_n13780 a_38716_n13780 0.012882f
C2203 a_27820_n16432 a_29161_n14476 0.042503f
C2204 a_47476_n14116 VDD 0.206217f
C2205 a_22820_n2804 a_25759_n3544 0.02738f
C2206 a_38403_n2367 a_38733_n2295 0.538085f
C2207 a_33292_n2716 a_33188_n2672 0.026665f
C2208 a_42660_n15304 a_42300_n15348 0.087066f
C2209 a_34248_n3310 a_34000_n3140 0.366988f
C2210 a_23844_n18440 VDD 0.208184f
C2211 a_44004_n16872 a_44092_n16916 0.285629f
C2212 a_44004_n4328 a_44092_n4372 0.285629f
C2213 OUT[2] OUT[3] 0.143354f
C2214 a_40060_n16916 a_40508_n16916 0.012882f
C2215 a_42076_n20485 VDD 0.329322f
C2216 a_37732_n18440 a_37372_n18484 0.087066f
C2217 a_26172_n18484 a_26060_n18917 0.026339f
C2218 a_45660_n5940 a_46108_n5940 0.012552f
C2219 a_27988_n4328 a_30871_n11728 0.401591f
C2220 a_39357_n5364 a_39500_n6373 0.031039f
C2221 a_47364_n5896 a_47452_n5940 0.285629f
C2222 a_27516_n20052 a_27964_n20052 0.012882f
C2223 a_28624_n9394 a_28644_n9815 0.484332f
C2224 a_29800_n9815 a_25724_n14564 0.181657f
C2225 a_27281_n16854 a_29992_n11150 0.032859f
C2226 a_46556_n9076 a_46668_n9509 0.026339f
C2227 a_27167_n10808 a_28121_n10980 0.014443f
C2228 a_28437_n13705 a_28009_n12168 0.024721f
C2229 a_45572_n9032 VDD 0.213324f
C2230 a_26635_n12996 a_26983_n12728 0.633318f
C2231 a_47812_n13736 a_47452_n13780 0.086635f
C2232 a_21772_n12996 a_21604_n15684 0.028863f
C2233 a_36588_n15348 VDD 0.321045f
C2234 a_47812_n15304 a_47900_n15348 0.285629f
C2235 a_46108_n15348 a_46556_n15348 0.012552f
C2236 a_31772_n18484 VDD 0.322689f
C2237 a_47452_n4372 a_47900_n4372 0.012001f
C2238 a_42436_n20388 VDD 0.203482f
C2239 a_33564_n18484 a_33452_n18917 0.026339f
C2240 a_44092_n18484 a_44540_n18484 0.012001f
C2241 a_34820_n20008 a_34460_n20052 0.087066f
C2242 a_39500_n7941 a_39860_n7844 0.086742f
C2243 a_46668_n7941 a_47116_n7941 0.012882f
C2244 a_40644_n2760 VDD 0.206914f
C2245 a_22220_n12996 a_25020_n11383 0.010114f
C2246 a_47004_n5940 VDD 0.313885f
C2247 a_39724_n11077 a_40172_n11077 0.012222f
C2248 a_41852_n20052 CLK 0.013107f
C2249 a_21892_n12952 VDD 0.820408f
C2250 a_22588_n2020 a_22918_n2020 0.75472f
C2251 a_21916_n1975 a_23954_n2020 0.03102f
C2252 a_47364_1944 OUT[5] 0.012298f
C2253 a_47452_n15348 VDD 0.313885f
C2254 a_25237_n4327 a_25759_n3544 0.471293f
C2255 a_23507_n2759 a_24233_n3980 0.016921f
C2256 a_25759_1944 a_25524_1243 0.061795f
C2257 a_35940_2475 a_36388_1944 0.206994f
C2258 a_21692_2431 a_22096_376 1.53613f
C2259 a_45572_n18440 VDD 0.213324f
C2260 a_37484_n17349 a_37932_n17349 0.012882f
C2261 a_44876_n6373 a_45324_n6373 0.012882f
C2262 a_37732_n20008 a_37820_n20052 0.285629f
C2263 a_41316_n20008 a_41764_n20008 0.013276f
C2264 a_28412_n20052 a_28300_n20485 0.026339f
C2265 a_26383_n2968 VDD 0.585754f
C2266 a_44428_n9509 a_44340_n9412 0.285629f
C2267 a_36500_n9412 a_36948_n9412 0.013276f
C2268 a_22220_n12996 a_28437_n13705 0.011689f
C2269 a_37859_377 VDD 1.5828f
C2270 a_46220_n6373 VDD 0.31977f
C2271 a_43084_n11077 a_42996_n10980 0.285629f
C2272 a_32158_n12212 a_33364_n11384 0.02303f
C2273 a_37844_n9412 VDD 0.214349f
C2274 a_45772_n12645 a_46220_n12645 0.012882f
C2275 a_26563_n12212 a_26532_n14437 0.01659f
C2276 a_24573_n12996 a_23816_n13248 0.032797f
C2277 a_36812_n12645 a_37172_n12548 0.087174f
C2278 a_47116_n12645 VDD 0.315469f
C2279 a_29295_n1400 a_29519_n1976 0.538085f
C2280 a_32413_n14564 a_33364_n14116 0.016516f
C2281 a_46668_n15781 VDD 0.318039f
C2282 a_45324_n15781 a_45772_n15781 0.012882f
C2283 a_34860_n3189 a_34552_n3140 0.934191f
C2284 a_30555_n2729 a_31787_n3969 0.052928f
C2285 a_37036_n15781 a_36948_n15684 0.285629f
C2286 a_42604_n2020 a_44764_n1669 0.012889f
C2287 a_22096_376 a_26284_1564 0.083445f
C2288 a_25524_1243 a_28153_1204 0.019043f
C2289 a_37484_n18917 VDD 0.322148f
C2290 a_25936_1564 a_26488_1564 0.361958f
C2291 a_27988_n20388 a_28324_n20008 0.011616f
C2292 a_23564_n20836 a_23844_n18820 0.036664f
C2293 a_38716_n4805 a_39164_n4805 0.012552f
C2294 a_37932_n17349 a_38292_n17252 0.087066f
C2295 a_22588_n18917 a_22948_n18820 0.087174f
C2296 a_36140_n18917 a_36588_n18917 0.012882f
C2297 a_37172_n7844 a_37284_n9032 0.026657f
C2298 a_24233_n8684 a_23816_n8544 0.633318f
C2299 a_22364_n8944 a_21872_n9394 0.011425f
C2300 a_44876_n3237 VDD 0.361572f
C2301 a_22264_n8988 a_22352_n12097 0.033982f
C2302 a_35064_1506 VDD 0.360568f
C2303 a_29476_n6980 VDD 0.591495f
C2304 a_45684_n10980 a_46132_n10980 0.013276f
C2305 a_28435_n10599 VDD 0.677206f
C2306 a_48012_n12645 a_47924_n12548 0.285629f
C2307 a_28752_n15348 a_27852_n14990 0.056398f
C2308 a_35156_n14116 a_35604_n14116 0.013276f
C2309 a_43980_n14213 a_43892_n14116 0.285629f
C2310 a_35940_n1931 a_36388_n1572 0.195342f
C2311 a_23844_n16872 VDD 0.211568f
C2312 a_26383_n2968 a_26271_n4306 0.033954f
C2313 a_43532_n3237 a_43980_n3237 0.012882f
C2314 a_47564_n15781 a_47924_n15684 0.087066f
C2315 a_34576_1204 a_34471_1575 0.536965f
C2316 a_33467_1116 a_34367_1619 0.116059f
C2317 a_31324_n4372 a_28492_332 0.020867f
C2318 a_32244_n18820 VDD 0.211974f
C2319 a_38292_n17252 a_38740_n17252 0.013276f
C2320 a_42324_n4 a_42157_n660 0.010897f
C2321 a_43980_n4805 a_43892_n4708 0.285629f
C2322 a_23479_n5156 a_21772_n9860 0.831259f
C2323 a_33900_n18917 a_33812_n18820 0.285629f
C2324 a_29308_n20485 a_29756_n20485 0.013103f
C2325 a_40956_n7508 VDD 0.330158f
C2326 a_39636_n10980 a_39524_n12168 0.026657f
C2327 a_24684_n16432 a_25559_n12548 0.021764f
C2328 a_38716_n10644 VDD 0.321613f
C2329 a_22016_n13665 a_22568_n13648 0.361958f
C2330 a_36140_n13780 VDD 0.296789f
C2331 a_43868_n1669 a_43780_n1572 0.285629f
C2332 a_38180_n16872 VDD 0.245127f
C2333 a_22500_n16872 a_22948_n16872 0.013276f
C2334 a_36052_n15684 a_36164_n16872 0.026657f
C2335 a_25636_n20008 VDD 0.210877f
C2336 a_42188_n6373 CLK 0.024601f
C2337 a_30900_n18820 a_31348_n18820 0.013276f
C2338 a_47924_n6276 a_47812_n7464 0.026657f
C2339 a_44428_n18917 a_44788_n18820 0.087066f
C2340 a_22264_n8988 a_21892_n9816 0.014899f
C2341 a_29756_n20485 a_29668_n20388 0.285629f
C2342 a_41316_n9032 a_41764_n9032 0.013276f
C2343 a_37732_n9032 a_37372_n9076 0.087066f
C2344 a_21872_n9394 a_22116_n9412 0.017382f
C2345 a_37680_n320 VDD 0.025442f
C2346 a_40956_n4372 VDD 0.330578f
C2347 a_47924_n9412 a_47812_n10600 0.026657f
C2348 a_30871_n11728 a_34652_n11391 0.016779f
C2349 a_35392_n10172 a_33900_n11428 0.212997f
C2350 a_37947_332 VDD 0.495014f
C2351 a_42636_n15781 CLK 0.01698f
C2352 a_36812_n7941 VDD 0.33038f
C2353 a_46132_n10980 a_46020_n12168 0.026657f
C2354 a_42548_n12548 a_42660_n13736 0.026657f
C2355 a_47004_n13780 VDD 0.313885f
C2356 a_27852_n14990 a_27316_n14820 0.393757f
C2357 a_24604_n17349 VDD 0.377558f
C2358 a_43444_n15684 a_43556_n16872 0.026657f
C2359 a_25600_n5895 a_25237_n5895 0.15208f
C2360 a_24913_864 a_25137_864 0.569174f
C2361 a_31772_n20052 VDD 0.337706f
C2362 a_27764_n18820 a_27876_n20008 0.026657f
C2363 a_39612_n7508 a_40060_n7508 0.012882f
C2364 a_43556_n7464 a_43644_n7508 0.285629f
C2365 a_23542_n1754 VDD 0.745127f
C2366 a_29668_n20388 a_30116_n20388 0.013276f
C2367 a_28617_n8548 a_25724_n14564 0.059092f
C2368 a_40732_n20485 a_41092_n20388 0.087174f
C2369 a_25020_n11383 a_28300_n15348 0.016844f
C2370 a_41316_n10600 a_41404_n10644 0.285629f
C2371 a_37372_n10644 a_37820_n10644 0.012882f
C2372 a_34576_1204 a_35156_n325 0.010214f
C2373 a_44788_n7844 VDD 0.22479f
C2374 a_39972_n12168 a_39612_n12212 0.087066f
C2375 a_36500_n10980 VDD 0.128512f
C2376 a_43725_908 a_43885_n452 0.018117f
C2377 a_22600_n12124 a_23564_n20836 0.056573f
C2378 a_34796_n13780 a_35244_n13780 0.012552f
C2379 a_21692_2431 a_26736_n364 0.05565f
C2380 a_42636_n14213 VDD 0.313885f
C2381 a_44228_n1572 a_44228_n2760 0.05841f
C2382 a_27988_n4328 a_29560_n3544 0.011718f
C2383 a_28436_n17252 VDD 0.203482f
C2384 a_36700_n16916 a_37284_n16872 0.016748f
C2385 a_43644_n705 a_43725_908 0.02964f
C2386 a_33533_908 a_34271_376 0.22442f
C2387 a_45572_n20008 VDD 0.213324f
C2388 a_40980_n5896 a_41068_n5940 0.285629f
C2389 a_34372_n18440 a_34012_n18484 0.087066f
C2390 a_34708_n18820 a_34820_n20008 0.026657f
C2391 a_24292_n20008 a_24740_n20008 0.013276f
C2392 a_37820_n7508 a_37708_n7941 0.026339f
C2393 a_42212_n10600 CLK 0.037136f
C2394 a_37632_n2020 VDD 0.468209f
C2395 a_21772_n9860 a_21892_n9816 0.389329f
C2396 a_22264_n8988 a_22568_n10512 0.049479f
C2397 a_24573_n9860 a_25642_n9816 0.014406f
C2398 a_24965_n9860 a_25237_n10599 0.018835f
C2399 a_38628_n4708 VDD 0.212303f
C2400 a_46916_n10600 a_46556_n10644 0.086742f
C2401 a_28437_n13705 a_28300_n15348 0.083583f
C2402 a_46020_n12168 a_46468_n12168 0.013276f
C2403 a_28009_n12168 VDD 0.500716f
C2404 a_42212_n13736 a_41852_n13780 0.087066f
C2405 a_34271_n1192 a_34895_n1192 0.104193f
C2406 a_47028_n14116 VDD 0.206217f
C2407 a_38268_n15348 a_38716_n15348 0.012882f
C2408 a_22820_n2804 a_25237_n4327 0.495937f
C2409 a_42212_n15304 a_42300_n15348 0.285629f
C2410 a_23396_n18440 VDD 0.209294f
C2411 a_44004_n16872 a_43644_n16916 0.087066f
C2412 a_31772_n16916 a_31660_n17349 0.026339f
C2413 a_44004_n4328 a_43644_n4372 0.086905f
C2414 a_39612_n4372 a_40060_n4372 0.013103f
C2415 a_41628_n20485 VDD 0.329322f
C2416 a_47364_n5896 a_47004_n5940 0.086742f
C2417 a_37284_n18440 a_37372_n18484 0.285629f
C2418 a_40868_n18440 a_41316_n18440 0.013276f
C2419 a_41652_n18820 a_41764_n20008 0.026657f
C2420 a_47004_n7508 a_47116_n7941 0.026339f
C2421 a_22164_n2760 VDD 0.953035f
C2422 a_27281_n16854 a_25724_n14564 0.041479f
C2423 a_44092_n10644 a_43980_n11077 0.026339f
C2424 a_27281_n16854 a_27639_n12537 0.048568f
C2425 a_45124_n9032 VDD 0.26277f
C2426 a_40508_n12212 a_40396_n12645 0.026339f
C2427 a_25573_n12167 a_25544_n16412 0.511924f
C2428 a_45660_n13780 a_46108_n13780 0.012552f
C2429 a_47364_n13736 a_47452_n13780 0.285629f
C2430 a_36140_n15348 VDD 0.296789f
C2431 a_42524_n2804 a_42972_n2804 0.013103f
C2432 a_47812_n15304 a_47452_n15348 0.086635f
C2433 a_24631_n3588 a_31348_n1931 0.111468f
C2434 a_31324_n18484 VDD 0.35151f
C2435 a_47452_n16916 a_47900_n16916 0.012001f
C2436 a_38716_n16916 a_38828_n17349 0.026339f
C2437 a_41988_n20388 VDD 0.203482f
C2438 a_45212_n5940 a_45324_n6373 0.026339f
C2439 a_34372_n20008 a_34460_n20052 0.285629f
C2440 a_30428_n20052 a_30876_n20052 0.012882f
C2441 a_39500_n7941 a_39412_n7844 0.285629f
C2442 a_39357_n2228 VDD 0.752706f
C2443 a_22264_n10556 a_22016_n10529 0.343433f
C2444 a_46556_n5940 VDD 0.31705f
C2445 a_22220_n12996 VDD 0.694653f
C2446 a_34572_n12645 a_35020_n12645 0.013103f
C2447 a_27744_n12908 VDD 1.85166f
C2448 a_21916_n1975 a_23542_n1754 0.034799f
C2449 a_33077_n1191 a_32308_n1976 0.025559f
C2450 a_29161_n14476 a_28752_n15348 0.129648f
C2451 a_47004_n15348 VDD 0.313885f
C2452 a_45660_n15348 a_45772_n15781 0.026339f
C2453 a_34348_n15781 a_34796_n15781 0.012882f
C2454 a_22164_n2760 a_26271_n4306 0.020796f
C2455 a_21692_2431 a_25936_1564 0.027008f
C2456 a_45124_n18440 VDD 0.26277f
C2457 a_47900_n16916 a_48012_n17349 0.026339f
C2458 a_40060_n18484 a_40172_n18917 0.026339f
C2459 a_43444_n7844 a_43892_n7844 0.013276f
C2460 a_37732_n20008 a_37372_n20052 0.087066f
C2461 a_43980_n9509 a_44340_n9412 0.087066f
C2462 a_45772_n6373 VDD 0.321879f
C2463 a_22220_n12996 a_21604_n13252 0.035085f
C2464 a_42636_n11077 a_42996_n10980 0.087066f
C2465 a_37396_n9412 VDD 0.211702f
C2466 a_36812_n12645 a_36724_n12548 0.285629f
C2467 a_46668_n12645 VDD 0.318039f
C2468 a_21772_n12996 a_25544_n16412 0.245388f
C2469 a_41292_n14213 a_41740_n14213 0.012882f
C2470 a_46220_n15781 VDD 0.31977f
C2471 a_36588_n15781 a_36948_n15684 0.087066f
C2472 a_34000_n3140 a_34552_n3140 0.361958f
C2473 a_47004_n2804 a_47116_n3237 0.026339f
C2474 a_42604_n2020 a_44316_n1669 0.012889f
C2475 a_25936_1564 a_26284_1564 0.401636f
C2476 a_25524_1243 a_27736_1248 0.042802f
C2477 a_37036_n18917 VDD 0.334604f
C2478 a_37932_n17349 a_37844_n17252 0.285629f
C2479 a_21792_n7464 a_21812_n6643 0.083468f
C2480 a_27988_n20388 a_27876_n20008 0.056574f
C2481 a_22588_n18917 a_22500_n18820 0.285629f
C2482 a_44788_n6276 a_45236_n6276 0.013276f
C2483 a_22876_n8988 a_21872_n9394 0.0189f
C2484 a_22016_n8961 a_24128_n8544 0.277491f
C2485 a_44092_n20052 a_44540_n20052 0.012001f
C2486 a_35356_n20052 a_35356_n20485 0.05841f
C2487 a_44428_n3237 VDD 0.323614f
C2488 a_34471_1575 VDD 0.798592f
C2489 a_47028_n9412 a_47476_n9412 0.013276f
C2490 a_47564_n12645 a_47924_n12548 0.087066f
C2491 a_38516_n12548 a_38964_n12548 0.013276f
C2492 a_22568_n13648 VDD 0.363142f
C2493 a_28752_n15348 a_27404_n14990 0.01003f
C2494 a_33077_n1191 a_34649_n2412 0.013139f
C2495 a_21916_n1975 a_22164_n2760 0.103642f
C2496 a_43532_n14213 a_43892_n14116 0.087066f
C2497 a_23396_n16872 VDD 0.210974f
C2498 a_47564_n15781 a_47476_n15684 0.285629f
C2499 a_38740_n15684 a_39188_n15684 0.013276f
C2500 a_33815_1384 a_34471_1575 0.510371f
C2501 a_28736_1944 a_28132_376 0.044473f
C2502 a_31796_n18820 VDD 0.21496f
C2503 a_43532_n4805 a_43892_n4708 0.087066f
C2504 a_46668_n18917 a_47116_n18917 0.012882f
C2505 a_33452_n18917 a_33812_n18820 0.087066f
C2506 a_25817_804 VDD 0.694495f
C2507 a_40508_n7508 VDD 0.315469f
C2508 a_38268_n10644 VDD 0.356786f
C2509 a_21604_n13252 a_22568_n13648 0.08126f
C2510 a_22016_n13665 a_22364_n13648 0.401636f
C2511 a_35692_n13780 VDD 0.296789f
C2512 a_43420_n1669 a_43780_n1572 0.087174f
C2513 a_45684_n14116 a_46132_n14116 0.013276f
C2514 a_37732_n16872 VDD 0.213126f
C2515 a_45236_n3140 a_45684_n3140 0.013276f
C2516 a_25188_n20008 VDD 0.215785f
C2517 a_42168_1564 a_42372_1564 0.66083f
C2518 a_32468_n17252 a_32580_n18440 0.026657f
C2519 a_24492_n5156 a_23949_n6724 0.02059f
C2520 a_24672_n11339 a_21812_n6643 0.079759f
C2521 a_22052_n18440 a_22500_n18440 0.013276f
C2522 a_41740_n6373 CLK 0.015046f
C2523 a_44428_n18917 a_44340_n18820 0.285629f
C2524 a_25612_n6679 a_29532_n10311 0.013551f
C2525 a_35119_n1170 VDD 0.325278f
C2526 a_37284_n9032 a_37372_n9076 0.285629f
C2527 a_23816_n8544 a_24573_n9860 0.022382f
C2528 a_29308_n20485 a_29668_n20388 0.087174f
C2529 a_37785_n364 VDD 0.502884f
C2530 a_42636_n12645 CLK 0.01698f
C2531 a_40508_n4372 VDD 0.296789f
C2532 a_33672_n10112 a_33900_n11428 0.03302f
C2533 a_35392_n10172 a_34652_n11391 0.55336f
C2534 a_36364_n7941 VDD 0.326475f
C2535 a_42188_n15781 CLK 0.047331f
C2536 a_30159_n13296 a_30555_n13780 0.018088f
C2537 a_46556_n13780 VDD 0.31705f
C2538 a_32860_n2020 a_37452_n3888 0.475368f
C2539 a_27404_n14990 a_27316_n14820 0.506857f
C2540 a_40532_n14116 a_40420_n15304 0.026657f
C2541 a_35156_n325 VDD 1.90627f
C2542 a_32580_n16872 a_33028_n16872 0.013276f
C2543 a_25600_n5895 a_24672_n11339 0.26228f
C2544 a_41204_n3140 a_41316_n4328 0.026657f
C2545 a_31324_n20052 VDD 0.368509f
C2546 a_39636_n17252 a_39524_n18440 0.026657f
C2547 a_43556_n7464 a_43196_n7508 0.087066f
C2548 a_41652_n18820 a_42100_n18820 0.013276f
C2549 a_22918_n2020 VDD 0.579732f
C2550 a_43644_n9076 a_44092_n9076 0.012882f
C2551 a_40732_n20485 a_40644_n20388 0.285629f
C2552 a_25831_n11428 a_27526_n9816 0.251728f
C2553 a_24180_n5112 VDD 0.894739f
C2554 a_41316_n10600 a_40956_n10644 0.087066f
C2555 a_28927_n10160 a_29332_n11301 0.010439f
C2556 a_44340_n7844 VDD 0.212126f
C2557 a_26563_n12212 a_27639_n12537 0.011052f
C2558 a_39524_n12168 a_39612_n12212 0.285629f
C2559 a_43556_n12168 a_44004_n12168 0.013276f
C2560 a_28300_n15348 VDD 1.20145f
C2561 a_21772_n12996 a_22140_n15348 0.011058f
C2562 a_22568_n1104 a_22772_n1104 0.66083f
C2563 a_22600_n12124 a_22948_n15684 0.017354f
C2564 a_36500_n13736 a_36588_n13780 0.285629f
C2565 a_42188_n14213 VDD 0.313885f
C2566 a_34796_n15348 a_35244_n15348 0.013103f
C2567 a_28454_n2424 a_27628_n3841 0.015853f
C2568 a_47476_n14116 a_47364_n15304 0.026657f
C2569 a_27988_n17252 VDD 0.11868f
C2570 a_47924_n3140 a_47812_n4328 0.026657f
C2571 a_33608_n4284 a_33416_n4240 0.934191f
C2572 a_45124_n20008 VDD 0.26277f
C2573 a_46580_n17252 a_46468_n18440 0.026657f
C2574 a_29980_n18484 a_30428_n18484 0.012882f
C2575 a_22444_n5156 a_33497_n9032 0.052446f
C2576 a_33924_n18440 a_34012_n18484 0.285629f
C2577 a_40980_n5896 a_40620_n5940 0.087174f
C2578 a_47004_n7508 a_47452_n7508 0.012222f
C2579 a_36388_n1572 VDD 0.647802f
C2580 a_40644_n20388 a_41092_n20388 0.013276f
C2581 a_22264_n8988 a_22364_n10512 0.015066f
C2582 a_38180_n4708 VDD 0.207244f
C2583 a_46468_n10600 a_46556_n10644 0.285629f
C2584 a_41764_n13736 a_41852_n13780 0.285629f
C2585 a_30408_n1104 a_30612_n1104 0.66083f
C2586 a_37820_n13780 a_38268_n13780 0.012882f
C2587 a_30159_n13296 a_31459_n14564 0.21163f
C2588 a_46580_n14116 VDD 0.209016f
C2589 a_42212_n15304 a_41852_n15348 0.087066f
C2590 a_22948_n18440 VDD 0.205626f
C2591 a_43556_n4328 a_43644_n4372 0.285629f
C2592 a_39612_n16916 a_40060_n16916 0.012882f
C2593 a_43556_n16872 a_43644_n16916 0.285629f
C2594 a_41180_n20485 VDD 0.329322f
C2595 a_45212_n5940 a_45660_n5940 0.012552f
C2596 a_46916_n5896 a_47004_n5940 0.285629f
C2597 a_25724_n18484 a_25612_n18917 0.026339f
C2598 a_27068_n20052 a_27516_n20052 0.012882f
C2599 a_21716_n2229 VDD 0.508071f
C2600 a_28617_n8548 a_30136_n10600 0.011663f
C2601 a_46108_n9076 a_46220_n9509 0.026339f
C2602 a_44540_n9076 VDD 0.353322f
C2603 a_26239_n12996 a_26635_n12996 0.025767f
C2604 a_44452_n12168 VDD 0.219497f
C2605 a_44228_n1192 a_44316_n1236 0.285629f
C2606 a_47364_n13736 a_47004_n13780 0.086742f
C2607 a_35692_n15348 VDD 0.296789f
C2608 a_47364_n15304 a_47452_n15348 0.285629f
C2609 a_45660_n15348 a_46108_n15348 0.012552f
C2610 a_24631_n3588 a_27988_n4328 0.255233f
C2611 a_30876_n18484 VDD 0.321966f
C2612 a_47004_n4372 a_47452_n4372 0.012222f
C2613 a_41540_n20388 VDD 0.203482f
C2614 a_43644_n18484 a_44092_n18484 0.012882f
C2615 a_46220_n7941 a_46668_n7941 0.012882f
C2616 a_39052_n7941 a_39412_n7844 0.087174f
C2617 a_34372_n20008 a_34012_n20052 0.087066f
C2618 a_38733_n2295 VDD 0.602387f
C2619 a_22264_n10556 a_21604_n10116 0.099099f
C2620 a_46108_n5940 VDD 0.318654f
C2621 a_39276_n11077 a_39724_n11077 0.013103f
C2622 a_29180_n9387 VDD 0.011991f
C2623 a_26983_n12728 VDD 1.32757f
C2624 a_21772_n12996 a_23564_n17700 0.232755f
C2625 a_28744_n14432 a_28752_n15348 0.032309f
C2626 a_21916_n1975 a_22918_n2020 0.024831f
C2627 a_34895_n1192 a_35288_n1975 0.010366f
C2628 a_44004_n1192 OUT[5] 0.073996f
C2629 a_46556_n15348 VDD 0.31705f
C2630 a_22164_n2760 a_26047_n4328 0.025161f
C2631 a_44540_n18484 VDD 0.353322f
C2632 a_37036_n17349 a_37484_n17349 0.012882f
C2633 a_44540_n4372 a_44428_n4805 0.026339f
C2634 a_44428_n6373 a_44876_n6373 0.012882f
C2635 a_39500_n6373 a_39412_n6276 0.285629f
C2636 a_40868_n20008 a_41316_n20008 0.013276f
C2637 a_37284_n20008 a_37372_n20052 0.285629f
C2638 a_25759_n3544 VDD 0.730699f
C2639 a_29800_n9815 a_29444_n10116 0.016045f
C2640 a_43980_n9509 a_43892_n9412 0.285629f
C2641 a_36388_1944 VDD 1.02237f
C2642 a_42548_n14116 CLK 0.029747f
C2643 a_45324_n6373 VDD 0.324845f
C2644 a_42636_n11077 a_42548_n10980 0.285629f
C2645 a_28121_n10980 a_27279_n12146 0.039161f
C2646 a_36948_n9412 VDD 0.21223f
C2647 a_45324_n12645 a_45772_n12645 0.012882f
C2648 a_36364_n12645 a_36724_n12548 0.087174f
C2649 a_46220_n12645 VDD 0.31977f
C2650 a_21772_n12996 a_23932_n16916 0.0107f
C2651 a_45772_n15781 VDD 0.321879f
C2652 a_44876_n15781 a_45324_n15781 0.012882f
C2653 a_36588_n15781 a_36500_n15684 0.285629f
C2654 a_34000_n3140 a_34348_n3140 0.401636f
C2655 a_24631_n3588 a_27628_n3841 0.218725f
C2656 a_42604_n2020 a_43868_n1669 0.01307f
C2657 a_36588_n18917 VDD 0.316762f
C2658 a_35940_2475 a_34576_1204 0.032681f
C2659 a_25936_1564 a_26796_1515 0.882105f
C2660 a_38268_n4805 a_38716_n4805 0.012552f
C2661 a_37484_n17349 a_37844_n17252 0.087066f
C2662 a_21792_n7464 a_22016_n6276 0.011348f
C2663 a_27988_n20388 a_27428_n20008 0.012624f
C2664 a_22140_n18917 a_22500_n18820 0.087174f
C2665 a_35692_n18917 a_36140_n18917 0.012882f
C2666 a_23564_n8292 a_23619_n9860 0.063042f
C2667 a_22264_n8988 a_21872_n9394 0.189518f
C2668 a_43980_n3237 VDD 0.32102f
C2669 a_25020_n11383 a_28927_n10160 0.030052f
C2670 a_28335_n10644 a_28435_n10599 0.264272f
C2671 a_45236_n10980 a_45684_n10980 0.013276f
C2672 a_42772_n4 a_42948_n1976 0.02146f
C2673 a_44004_n1192 a_42948_n1976 0.056916f
C2674 a_47564_n12645 a_47476_n12548 0.285629f
C2675 a_22364_n13648 VDD 0.010384f
C2676 a_34708_n14116 a_35156_n14116 0.013276f
C2677 a_43532_n14213 a_43444_n14116 0.285629f
C2678 a_27820_n16432 a_27709_n16132 0.066658f
C2679 a_21916_n1975 a_21716_n2229 0.015226f
C2680 a_22948_n16872 VDD 0.205195f
C2681 a_47116_n15781 a_47476_n15684 0.087066f
C2682 a_43084_n3237 a_43532_n3237 0.012882f
C2683 a_28736_1944 a_28492_332 0.029938f
C2684 a_22500_n1976 a_28132_376 0.042033f
C2685 a_33467_1116 a_34471_1575 0.020455f
C2686 a_31348_n18820 VDD 0.239843f
C2687 a_37844_n17252 a_38292_n17252 0.013276f
C2688 a_43532_n4805 a_43444_n4708 0.285629f
C2689 a_33452_n18917 a_33364_n18820 0.285629f
C2690 a_40308_n6276 a_40420_n7464 0.026657f
C2691 a_25573_n12167 a_25831_n11428 0.478254f
C2692 a_47452_1900 EOC 0.024173f
C2693 a_22772_n4240 VDD 0.299834f
C2694 a_27485_n10068 a_28247_n10599 0.045583f
C2695 a_28437_n13705 a_28927_n10160 0.227134f
C2696 a_40532_n9412 a_40420_n10600 0.026657f
C2697 a_25137_864 VDD 0.256813f
C2698 a_40060_n7508 VDD 0.316003f
C2699 a_39188_n10980 a_39076_n12168 0.026657f
C2700 a_24965_n9860 a_25636_n14520 0.581944f
C2701 a_26736_n364 a_26631_7 0.536965f
C2702 a_37820_n10644 VDD 0.322978f
C2703 a_22016_n13665 a_22876_n13692 0.882105f
C2704 a_21604_n13252 a_22364_n13648 0.011851f
C2705 a_35244_n13780 VDD 0.296789f
C2706 a_43420_n1669 a_43332_n1572 0.285629f
C2707 a_31324_n4372 a_31968_n704 0.010829f
C2708 a_37284_n16872 VDD 0.231657f
C2709 a_22052_n16872 a_22500_n16872 0.013276f
C2710 a_35604_n15684 a_35716_n16872 0.026657f
C2711 a_42476_1515 a_43416_1248 0.056721f
C2712 a_41616_1564 a_43728_1248 0.277491f
C2713 a_24740_n20008 VDD 0.235926f
C2714 a_23887_n5156 a_23949_n6724 0.024936f
C2715 a_41292_n6373 CLK 0.01454f
C2716 a_30452_n18820 a_30900_n18820 0.013276f
C2717 a_43980_n18917 a_44340_n18820 0.087066f
C2718 a_47476_n6276 a_47364_n7464 0.026657f
C2719 a_34895_n1192 VDD 0.582344f
C2720 a_40868_n9032 a_41316_n9032 0.013276f
C2721 a_29308_n20485 a_29220_n20388 0.285629f
C2722 a_37368_n320 VDD 1.36854f
C2723 a_40060_n4372 VDD 0.297323f
C2724 a_42188_n12645 CLK 0.047331f
C2725 a_25020_n11383 a_29332_n11301 0.027797f
C2726 a_47476_n9412 a_47364_n10600 0.026657f
C2727 a_30104_n1148 VDD 0.842001f
C2728 a_33672_n10112 a_34652_n11391 0.07946f
C2729 a_34089_n10252 a_33900_n11428 0.013432f
C2730 a_45684_n10980 a_45572_n12168 0.026657f
C2731 a_36612_n12168 a_36700_n12212 0.285629f
C2732 a_42100_n12548 a_42212_n13736 0.026657f
C2733 a_46108_n13780 VDD 0.318654f
C2734 a_28752_n15348 a_28568_n16066 0.612085f
C2735 a_47900_n16916 VDD 0.335152f
C2736 a_42996_n15684 a_43108_n16872 0.026657f
C2737 a_30876_n20052 VDD 0.336983f
C2738 a_25724_n18484 a_26172_n18484 0.012001f
C2739 a_39164_n7508 a_39612_n7508 0.012882f
C2740 a_33497_n9032 a_33308_n7376 0.03f
C2741 a_43108_n7464 a_43196_n7508 0.285629f
C2742 a_21812_n6643 a_25860_n9032 0.049741f
C2743 a_27316_n18820 a_27428_n20008 0.026657f
C2744 a_40060_n20485 a_40644_n20388 0.016748f
C2745 a_29220_n20388 a_29668_n20388 0.013276f
C2746 a_25831_n11428 a_27302_n9816 0.035528f
C2747 a_25724_n14564 a_24152_n11680 0.016041f
C2748 a_40868_n10600 a_40956_n10644 0.285629f
C2749 a_43892_n7844 VDD 0.210071f
C2750 a_39524_n12168 a_39164_n12212 0.087066f
C2751 a_23564_n11428 a_24128_n13248 0.04547f
C2752 a_34538_n10980 VDD 0.014549f
C2753 a_22600_n12124 a_22500_n15684 0.056315f
C2754 a_21772_n12996 a_21692_n15348 0.047171f
C2755 a_36500_n13736 a_36140_n13780 0.086635f
C2756 a_41740_n14213 VDD 0.313885f
C2757 a_43780_n1572 a_43780_n2760 0.05841f
C2758 a_24516_n17252 VDD 0.242179f
C2759 a_33015_n4284 a_33416_n4240 0.882105f
C2760 a_36252_n16916 a_36700_n16916 0.012001f
C2761 a_44540_n20052 VDD 0.334642f
C2762 a_43668_n5896 a_44116_n5896 0.013276f
C2763 a_33924_n18440 a_33564_n18484 0.087066f
C2764 a_40532_n5896 a_40620_n5940 0.285629f
C2765 a_23844_n20008 a_24292_n20008 0.013276f
C2766 a_34260_n18820 a_34372_n20008 0.026657f
C2767 a_37372_n7508 a_37260_n7941 0.026339f
C2768 a_36744_n1954 VDD 0.652815f
C2769 a_24573_n9860 a_24965_n9860 0.464885f
C2770 a_46468_n10600 a_46108_n10644 0.086905f
C2771 a_45572_n12168 a_46020_n12168 0.013276f
C2772 a_41764_n13736 a_41404_n13780 0.087066f
C2773 a_46132_n14116 VDD 0.210512f
C2774 a_41764_n15304 a_41852_n15348 0.285629f
C2775 a_37820_n15348 a_38268_n15348 0.012882f
C2776 a_31392_n2760 a_31636_n2760 0.015253f
C2777 a_22500_n1976 a_23507_n2759 0.455099f
C2778 a_22500_n18440 VDD 0.203482f
C2779 a_31324_n16916 a_31212_n17349 0.026339f
C2780 a_39164_n4372 a_39612_n4372 0.013103f
C2781 a_43556_n16872 a_43196_n16916 0.087066f
C2782 a_43556_n4328 a_43196_n4372 0.086905f
C2783 a_40732_n20485 VDD 0.333995f
C2784 a_46916_n5896 a_46556_n5940 0.086742f
C2785 a_40420_n18440 a_40868_n18440 0.013276f
C2786 a_46556_n7508 a_46668_n7941 0.026339f
C2787 a_41204_n18820 a_41316_n20008 0.026657f
C2788 a_31341_n8292 a_31965_n8292 0.104193f
C2789 a_22820_n2804 VDD 1.46259f
C2790 a_43644_n10644 a_43532_n11077 0.026339f
C2791 a_35816_n174 a_35156_n325 0.10802f
C2792 a_42948_n1976 a_42244_n1572 0.226094f
C2793 a_44092_n9076 VDD 0.3211f
C2794 a_40060_n12212 a_39948_n12645 0.026339f
C2795 a_44004_n12168 VDD 0.2108f
C2796 a_24684_n16432 a_24604_n17349 0.02963f
C2797 a_46916_n13736 a_47004_n13780 0.285629f
C2798 a_45212_n13780 a_45660_n13780 0.012552f
C2799 a_35244_n15348 VDD 0.296789f
C2800 a_47364_n15304 a_47004_n15348 0.086742f
C2801 a_42076_n2804 a_42524_n2804 0.013103f
C2802 a_40652_n1572 a_45660_n1669 0.019548f
C2803 a_30428_n18484 VDD 0.319233f
C2804 a_47004_n16916 a_47452_n16916 0.012222f
C2805 a_38268_n16916 a_38380_n17349 0.026339f
C2806 a_41092_n20388 VDD 0.203482f
C2807 a_32668_n18484 a_32780_n18917 0.026339f
C2808 a_29980_n20052 a_30428_n20052 0.012882f
C2809 a_33924_n20008 a_34012_n20052 0.285629f
C2810 a_39052_n7941 a_38964_n7844 0.285629f
C2811 a_38403_n2367 VDD 0.358606f
C2812 a_22220_n12996 a_28335_n10644 0.704419f
C2813 a_40172_n9509 a_40620_n9509 0.012222f
C2814 a_23479_n5156 a_27192_n14286 0.156737f
C2815 a_45660_n5940 VDD 0.320877f
C2816 a_28868_n9387 VDD 0.021926f
C2817 a_34124_n12645 a_34572_n12645 0.013103f
C2818 a_26635_n12996 VDD 0.464719f
C2819 a_21828_n1931 a_22588_n2020 0.010062f
C2820 a_46108_n15348 VDD 0.318654f
C2821 a_33900_n15781 a_34348_n15781 0.012882f
C2822 a_45212_n15348 a_45324_n15781 0.026339f
C2823 a_22164_n2760 a_25423_n4328 0.031572f
C2824 a_44092_n18484 VDD 0.3211f
C2825 a_24836_n4708 a_24180_n5112 0.015646f
C2826 a_47452_n16916 a_47564_n17349 0.026339f
C2827 a_39612_n18484 a_39724_n18917 0.026339f
C2828 a_24380_n18917 a_24828_n18917 0.013103f
C2829 a_21812_n6643 a_22712_n7420 0.0455f
C2830 a_42996_n7844 a_43444_n7844 0.013276f
C2831 a_25237_n4327 VDD 1.53085f
C2832 a_27281_n16854 a_29444_n10116 0.044865f
C2833 a_43532_n9509 a_43892_n9412 0.087066f
C2834 a_35940_2475 VDD 0.485509f
C2835 a_42100_n14116 CLK 0.020589f
C2836 a_44876_n6373 VDD 0.360805f
C2837 a_42188_n11077 a_42548_n10980 0.087066f
C2838 a_36500_n9412 VDD 0.129651f
C2839 a_36364_n12645 a_36276_n12548 0.285629f
C2840 a_23564_n11428 a_24220_n15260 0.011215f
C2841 a_45772_n12645 VDD 0.321879f
C2842 a_21772_n12996 a_23484_n16916 0.014859f
C2843 a_45324_n15781 VDD 0.324845f
C2844 a_46556_n2804 a_46668_n3237 0.026339f
C2845 a_36140_n15781 a_36500_n15684 0.087066f
C2846 a_34000_n3140 a_34860_n3189 0.882105f
C2847 a_42604_n2020 a_43420_n1669 0.013252f
C2848 a_25524_1243 a_26488_1564 0.08126f
C2849 a_36140_n18917 VDD 0.313885f
C2850 a_25936_1564 a_22096_376 0.337386f
C2851 a_47564_n17349 a_48012_n17349 0.012882f
C2852 a_37484_n17349 a_37396_n17252 0.285629f
C2853 a_44340_n6276 a_44788_n6276 0.013276f
C2854 a_22140_n18917 a_22052_n18820 0.285629f
C2855 a_43644_n20052 a_44092_n20052 0.012882f
C2856 a_34908_n20052 a_34908_n20485 0.05841f
C2857 a_23564_n8292 a_21772_n9860 0.014374f
C2858 a_22016_n8961 a_21872_n9394 0.064587f
C2859 a_43532_n3237 VDD 0.319276f
C2860 a_25020_n11383 a_28437_n13705 0.031782f
C2861 a_46580_n9412 a_47028_n9412 0.013276f
C2862 a_23220_n7376 VDD 0.300454f
C2863 a_28927_n10160 VDD 1.20198f
C2864 a_44004_n1192 a_44509_n452 0.013272f
C2865 a_38068_n12548 a_38516_n12548 0.013276f
C2866 a_47116_n12645 a_47476_n12548 0.087066f
C2867 a_22876_n13692 VDD 0.248837f
C2868 a_43084_n14213 a_43444_n14116 0.087066f
C2869 a_21916_n1975 a_22820_n2804 0.199727f
C2870 a_35288_n1975 a_35940_n1931 0.114265f
C2871 a_22500_n16872 VDD 0.203482f
C2872 a_25237_n4327 a_26271_n4306 0.057826f
C2873 a_38292_n15684 a_38740_n15684 0.013276f
C2874 a_47116_n15781 a_47028_n15684 0.285629f
C2875 a_22500_n1976 a_28492_332 0.113276f
C2876 a_30900_n18820 VDD 0.2134f
C2877 a_43084_n4805 a_43444_n4708 0.087066f
C2878 a_46220_n18917 a_46668_n18917 0.012882f
C2879 a_27988_n4328 a_30787_n12167 0.129753f
C2880 a_32780_n18917 a_33364_n18820 0.016748f
C2881 a_28617_n8548 a_28225_n9031 0.270381f
C2882 a_47364_1944 EOC 0.049294f
C2883 a_24128_n3840 VDD 0.024681f
C2884 a_24913_864 VDD 0.297901f
C2885 a_39612_n7508 VDD 0.31906f
C2886 a_27279_n12146 a_28009_n12168 0.212426f
C2887 a_24964_n14116 a_28040_n12493 0.016098f
C2888 a_25975_n184 a_26631_7 0.510371f
C2889 a_37372_n10644 VDD 0.327457f
C2890 a_21604_n13252 a_22876_n13692 0.05539f
C2891 a_34796_n13780 VDD 0.300786f
C2892 a_42244_n1572 a_43332_n1572 0.016177f
C2893 a_45236_n14116 a_45684_n14116 0.013276f
C2894 a_36700_n16916 VDD 0.347096f
C2895 a_44788_n3140 a_45236_n3140 0.013276f
C2896 a_42476_1515 a_42372_1564 0.026665f
C2897 a_41616_1564 a_43833_1204 0.020455f
C2898 a_24292_n20008 VDD 0.212186f
C2899 a_41964_1564 a_42168_1564 0.048436f
C2900 a_21604_n18440 a_22052_n18440 0.013276f
C2901 a_32020_n17252 a_32132_n18440 0.026657f
C2902 a_40396_n6373 CLK 0.014423f
C2903 a_43980_n18917 a_43892_n18820 0.285629f
C2904 a_34271_n1192 VDD 0.72072f
C2905 a_39612_n20485 a_40060_n20485 0.013103f
C2906 a_39612_n4372 VDD 0.30038f
C2907 a_25020_n11383 a_27391_n11384 0.028633f
C2908 a_34089_n10252 a_34652_n11391 0.19022f
C2909 a_31965_n8292 VDD 0.713343f
C2910 a_36612_n12168 a_36252_n12212 0.086905f
C2911 a_29332_n11301 VDD 1.86087f
C2912 a_45660_n13780 VDD 0.320877f
C2913 a_40084_n14116 a_39972_n15304 0.026657f
C2914 a_47452_n16916 VDD 0.313885f
C2915 a_32132_n16872 a_32580_n16872 0.013276f
C2916 a_30428_n20052 VDD 0.33425f
C2917 a_39188_n17252 a_39076_n18440 0.026657f
C2918 a_41204_n18820 a_41652_n18820 0.013276f
C2919 a_21812_n6643 a_25412_n8501 0.491366f
C2920 a_43108_n7464 a_42748_n7508 0.087066f
C2921 a_22588_n2020 VDD 0.307292f
C2922 a_40060_n20485 a_39972_n20388 0.285629f
C2923 a_43196_n9076 a_43644_n9076 0.012882f
C2924 a_25724_n14564 a_24569_n11820 0.042768f
C2925 a_40868_n10600 a_40508_n10644 0.087066f
C2926 a_43444_n7844 VDD 0.208665f
C2927 a_43108_n12168 a_43556_n12168 0.013276f
C2928 a_27279_n12146 a_27744_n12908 0.021762f
C2929 a_39076_n12168 a_39164_n12212 0.285629f
C2930 a_25880_n11708 a_25831_n12996 0.015514f
C2931 a_44004_n1192 a_43555_n452 0.072896f
C2932 a_36052_n13736 a_36140_n13780 0.285629f
C2933 a_22600_n12124 a_22052_n15684 0.013246f
C2934 a_22876_n1148 a_22772_n1104 0.026665f
C2935 a_41292_n14213 VDD 0.318502f
C2936 a_34348_n15348 a_34796_n15348 0.013103f
C2937 a_47028_n14116 a_46916_n15304 0.026657f
C2938 a_48012_n17349 VDD 0.343411f
C2939 a_47476_n3140 a_47364_n4328 0.026657f
C2940 a_33120_n3884 a_33416_n4240 0.05539f
C2941 a_32909_841 a_33533_908 0.104193f
C2942 a_44092_n20052 VDD 0.335452f
C2943 a_26631_7 a_27032_51 0.882105f
C2944 a_33476_n18440 a_33564_n18484 0.285629f
C2945 a_29532_n18484 a_29980_n18484 0.012882f
C2946 a_46132_n17252 a_46020_n18440 0.026657f
C2947 a_40532_n5896 a_40172_n5940 0.087174f
C2948 a_46556_n7508 a_47004_n7508 0.012222f
C2949 a_35940_n1931 VDD 0.460335f
C2950 a_23949_n9860 a_24965_n9860 0.082276f
C2951 a_22264_n8988 a_22016_n10529 0.03054f
C2952 a_47364_n10600 a_47812_n10600 0.013276f
C2953 a_46020_n10600 a_46108_n10644 0.285629f
C2954 a_25880_n11708 VDD 0.447309f
C2955 a_37372_n13780 a_37820_n13780 0.012882f
C2956 a_41316_n13736 a_41404_n13780 0.285629f
C2957 a_30716_n1148 a_30612_n1104 0.026665f
C2958 a_45684_n14116 VDD 0.212747f
C2959 a_37221_n3543 a_37585_n3140 0.019999f
C2960 a_31412_n2276 a_31636_n2760 0.013419f
C2961 a_41764_n15304 a_41404_n15348 0.087066f
C2962 a_22052_n18440 VDD 0.203482f
C2963 a_43108_n16872 a_43196_n16916 0.285629f
C2964 a_39164_n16916 a_39612_n16916 0.012882f
C2965 a_43108_n4328 a_43196_n4372 0.285629f
C2966 a_35816_n174 a_30104_n1148 0.024556f
C2967 a_40060_n20485 VDD 0.325703f
C2968 a_46468_n5896 a_46556_n5940 0.285629f
C2969 a_26620_n20052 a_27068_n20052 0.012882f
C2970 a_30676_n7844 a_31965_n8292 0.024857f
C2971 a_45660_n9076 a_45772_n9509 0.026339f
C2972 a_27526_n9816 a_25724_n14564 0.020901f
C2973 a_28624_n9394 a_22220_n12996 0.088593f
C2974 a_36773_n5468 VDD 0.74365f
C2975 a_43644_n9076 VDD 0.319164f
C2976 a_25831_n12996 a_26239_n12996 0.070482f
C2977 a_43556_n12168 VDD 0.209225f
C2978 a_46916_n13736 a_46556_n13780 0.086742f
C2979 a_34796_n15348 VDD 0.296789f
C2980 a_46916_n15304 a_47004_n15348 0.285629f
C2981 a_45212_n15348 a_45660_n15348 0.012552f
C2982 a_40652_n1572 a_45212_n1669 0.033754f
C2983 a_24631_n3588 a_30584_n1954 0.037891f
C2984 a_26527_51 VDD 0.022335f
C2985 a_29980_n18484 VDD 0.317392f
C2986 a_46556_n4372 a_47004_n4372 0.012222f
C2987 a_22052_n4708 a_29612_n8292 0.035521f
C2988 a_40644_n20388 VDD 0.224235f
C2989 a_42324_n4 a_42772_n4 0.013276f
C2990 a_43196_n18484 a_43644_n18484 0.012882f
C2991 a_45772_n7941 a_46220_n7941 0.012882f
C2992 a_33924_n20008 a_33564_n20052 0.087066f
C2993 a_23564_n8292 a_22016_n8961 0.036036f
C2994 a_47924_n18820 a_47812_n20008 0.026657f
C2995 a_38604_n7941 a_38964_n7844 0.087174f
C2996 a_23479_n5156 a_26944_n14116 0.058721f
C2997 a_45212_n5940 VDD 0.344357f
C2998 a_38828_n11077 a_39276_n11077 0.013103f
C2999 a_26239_n12996 VDD 0.542695f
C3000 a_21916_n1975 a_22588_n2020 0.0644f
C3001 a_34271_n1192 a_34223_n1976 0.012956f
C3002 a_44540_n13780 a_44428_n14213 0.026339f
C3003 a_45660_n15348 VDD 0.320877f
C3004 a_22164_n2760 a_23816_n3840 0.035626f
C3005 a_43644_n18484 VDD 0.319164f
C3006 a_21692_2431 a_25524_1243 0.01894f
C3007 a_36588_n17349 a_37036_n17349 0.012882f
C3008 a_44092_n4372 a_43980_n4805 0.026339f
C3009 a_22220_n9860 a_24180_n5112 0.41982f
C3010 a_21812_n6643 a_22464_n7393 0.024554f
C3011 a_43980_n6373 a_44428_n6373 0.012882f
C3012 a_40420_n20008 a_40868_n20008 0.013276f
C3013 a_35120_n9412 a_25020_n11383 0.024086f
C3014 a_25831_n11428 a_24964_n14116 0.427862f
C3015 a_43532_n9509 a_43444_n9412 0.285629f
C3016 a_44428_n6373 VDD 0.336571f
C3017 a_42188_n11077 a_42100_n10980 0.285629f
C3018 a_28437_n13705 a_25831_n12996 0.231611f
C3019 a_25020_n11383 VDD 0.94103f
C3020 a_44876_n12645 a_45324_n12645 0.012882f
C3021 a_23564_n11428 a_23608_n15260 0.165195f
C3022 a_35916_n12645 a_36276_n12548 0.087174f
C3023 a_45324_n12645 VDD 0.324845f
C3024 a_21772_n12996 a_23036_n16916 0.015944f
C3025 a_44876_n15781 VDD 0.360805f
C3026 a_44428_n15781 a_44876_n15781 0.012882f
C3027 a_36140_n15781 a_36052_n15684 0.285629f
C3028 a_24631_n3588 a_31292_n2804 0.216675f
C3029 a_42604_n2020 a_42244_n1572 0.58411f
C3030 a_25524_1243 a_26284_1564 0.011851f
C3031 a_35692_n18917 VDD 0.313885f
C3032 a_37036_n17349 a_37396_n17252 0.087066f
C3033 a_21692_n18917 a_22052_n18820 0.087174f
C3034 a_35244_n18917 a_35692_n18917 0.012882f
C3035 a_21604_n8548 a_21872_n9394 0.01586f
C3036 a_43084_n3237 VDD 0.315943f
C3037 a_34576_1204 VDD 1.80044f
C3038 a_24576_n6976 VDD 0.035526f
C3039 a_44788_n10980 a_45236_n10980 0.013276f
C3040 a_28437_n13705 VDD 0.702437f
C3041 a_44004_n1192 a_43885_n452 0.044043f
C3042 a_47116_n12645 a_47028_n12548 0.285629f
C3043 a_22016_n13665 VDD 0.808632f
C3044 a_43084_n14213 a_42996_n14116 0.285629f
C3045 a_34260_n14116 a_34708_n14116 0.013276f
C3046 a_22052_n16872 VDD 0.203482f
C3047 a_25237_n4327 a_26047_n4328 0.060003f
C3048 a_42636_n3237 a_43084_n3237 0.012882f
C3049 a_46668_n15781 a_47028_n15684 0.087066f
C3050 a_44004_n1192 a_43644_n705 0.347961f
C3051 a_33815_1384 a_34576_1204 0.042802f
C3052 a_30452_n18820 VDD 0.211196f
C3053 a_43084_n4805 a_42996_n4708 0.285629f
C3054 a_37396_n17252 a_37844_n17252 0.013276f
C3055 a_48012_n17349 a_47924_n17252 0.285629f
C3056 a_45236_n4 VDD 0.147845f
C3057 a_39860_n6276 a_39972_n7464 0.026657f
C3058 a_32780_n18917 a_32692_n18820 0.285629f
C3059 a_40084_n9412 a_39972_n10600 0.026657f
C3060 a_27281_n16854 a_28121_n10980 0.606898f
C3061 a_39164_n7508 VDD 0.320421f
C3062 a_27055_n12168 a_28009_n12168 0.014972f
C3063 a_38740_n10980 a_38628_n12168 0.026657f
C3064 a_25975_n184 a_26736_n364 0.042802f
C3065 a_25627_n452 a_26631_7 0.020455f
C3066 a_44452_n10600 VDD 0.219497f
C3067 a_21604_n13252 a_22016_n13665 0.536965f
C3068 a_22600_n12124 a_23608_n15260 0.018075f
C3069 a_33280_n13248 VDD 0.010444f
C3070 a_42244_n1572 a_42448_n1572 0.033243f
C3071 a_36252_n16916 VDD 0.315469f
C3072 a_35156_n15684 a_35268_n16872 0.026657f
C3073 a_21604_n16872 a_22052_n16872 0.013276f
C3074 a_41616_1564 a_43416_1248 0.510371f
C3075 a_42476_1515 a_42168_1564 0.934191f
C3076 a_23844_n20008 VDD 0.208184f
C3077 a_23887_n5156 a_21812_n6643 0.79627f
C3078 a_22544_n4690 a_24573_n6724 0.466048f
C3079 a_47476_n4708 a_47924_n4708 0.013276f
C3080 a_39948_n6373 CLK 0.014191f
C3081 a_30004_n18820 a_30452_n18820 0.013276f
C3082 a_47028_n6276 a_46916_n7464 0.026657f
C3083 a_43532_n18917 a_43892_n18820 0.087066f
C3084 a_33252_n1192 VDD 0.581644f
C3085 a_28300_n20485 a_28212_n20388 0.285629f
C3086 a_40420_n9032 a_40868_n9032 0.013276f
C3087 a_39164_n4372 VDD 0.307463f
C3088 a_25020_n11383 a_27167_n10808 0.029444f
C3089 a_47028_n9412 a_46916_n10600 0.026657f
C3090 a_31341_n8292 VDD 0.607655f
C3091 a_36164_n12168 a_36252_n12212 0.285629f
C3092 a_45236_n10980 a_45124_n12168 0.026657f
C3093 a_27391_n11384 VDD 0.326784f
C3094 a_41652_n12548 a_41764_n13736 0.026657f
C3095 a_45212_n13780 VDD 0.342281f
C3096 a_47004_n16916 VDD 0.313885f
C3097 a_27988_n4328 a_25612_n6679 0.029801f
C3098 a_40308_n3140 a_40420_n4328 0.026657f
C3099 a_42548_n15684 a_42660_n16872 0.026657f
C3100 a_29980_n20052 VDD 0.332409f
C3101 a_25276_n18484 a_25724_n18484 0.012222f
C3102 a_42660_n7464 a_42748_n7508 0.285629f
C3103 a_26868_n18820 a_26980_n20008 0.026657f
C3104 a_38716_n7508 a_39164_n7508 0.012882f
C3105 a_21828_n1931 VDD 0.489685f
C3106 a_25573_n12167 a_25724_n14564 1.51956f
C3107 a_39612_n20485 a_39972_n20388 0.087174f
C3108 a_22564_n5112 VDD 0.79393f
C3109 a_25020_n11383 a_32158_n12212 0.03956f
C3110 a_44004_n10600 a_44452_n10600 0.013276f
C3111 a_40420_n10600 a_40508_n10644 0.285629f
C3112 a_42996_n7844 VDD 0.205948f
C3113 a_39076_n12168 a_38716_n12212 0.087066f
C3114 a_42860_n101 a_42772_n4 0.285629f
C3115 a_36052_n13736 a_35692_n13780 0.086905f
C3116 a_21772_n12996 a_22052_n15304 0.014571f
C3117 a_40620_n14213 VDD 0.344269f
C3118 a_43332_n1572 a_43332_n2760 0.05841f
C3119 a_47564_n17349 VDD 0.315469f
C3120 a_35804_n16916 a_36252_n16916 0.012222f
C3121 a_33015_n4284 a_32911_n4240 0.277491f
C3122 a_43644_n20052 VDD 0.332597f
C3123 a_26736_n364 a_27032_51 0.05539f
C3124 a_28132_376 a_28336_376 0.033243f
C3125 a_33476_n18440 a_33116_n18484 0.087066f
C3126 a_43220_n5896 a_43668_n5896 0.013276f
C3127 a_40084_n5896 a_40172_n5940 0.285629f
C3128 a_22264_n5852 a_23949_n6724 0.013814f
C3129 a_42660_n7464 CLK 0.017841f
C3130 a_33812_n18820 a_33924_n20008 0.026657f
C3131 a_23396_n20008 a_23844_n20008 0.013276f
C3132 a_35288_n1975 VDD 0.454189f
C3133 a_23949_n9860 a_24573_n9860 0.104193f
C3134 a_22264_n8988 a_21604_n10116 0.016035f
C3135 a_33900_n11428 a_34350_n10980 0.011098f
C3136 a_46020_n10600 a_45660_n10644 0.086905f
C3137 a_32767_n9010 VDD 0.325642f
C3138 a_45124_n12168 a_45572_n12168 0.013276f
C3139 a_23108_n12080 VDD 0.300922f
C3140 a_41316_n13736 a_40956_n13780 0.087066f
C3141 a_45236_n14116 VDD 0.229781f
C3142 a_37221_n3543 a_22052_n4708 0.079637f
C3143 a_41316_n15304 a_41404_n15348 0.285629f
C3144 a_37372_n15348 a_37820_n15348 0.012882f
C3145 a_21604_n18440 VDD 0.223768f
C3146 a_43108_n16872 a_42748_n16916 0.087066f
C3147 a_43108_n4328 a_42748_n4372 0.086905f
C3148 a_30876_n16916 a_30764_n17349 0.026339f
C3149 a_39612_n20485 VDD 0.30038f
C3150 a_46468_n5896 a_46108_n5940 0.086905f
C3151 a_24828_n18484 a_24828_n18917 0.05841f
C3152 a_39972_n18440 a_40420_n18440 0.013276f
C3153 a_46108_n7508 a_46220_n7941 0.026339f
C3154 a_29800_n9815 a_22220_n12996 0.195671f
C3155 a_27302_n9816 a_25724_n14564 0.01308f
C3156 a_25573_n12167 a_25237_n13735 0.028241f
C3157 a_43196_n10644 a_43084_n11077 0.026339f
C3158 a_27167_n10808 a_27391_n11384 0.538085f
C3159 a_43196_n9076 VDD 0.316157f
C3160 a_39612_n12212 a_39500_n12645 0.026339f
C3161 a_43108_n12168 VDD 0.206217f
C3162 a_46468_n13736 a_46556_n13780 0.285629f
C3163 a_34348_n15348 VDD 0.296789f
C3164 a_46916_n15304 a_46556_n15348 0.086742f
C3165 a_41628_n2804 a_42076_n2804 0.013103f
C3166 a_40652_n1572 a_44764_n1669 0.019181f
C3167 a_27224_n62 VDD 0.360568f
C3168 a_29532_n18484 VDD 0.320804f
C3169 a_46556_n16916 a_47004_n16916 0.012222f
C3170 a_37820_n16916 a_37932_n17349 0.026339f
C3171 a_39972_n20388 VDD 0.211023f
C3172 a_25612_n6679 a_29123_n6679 0.037813f
C3173 a_32220_n18484 a_32332_n18917 0.026339f
C3174 a_38604_n7941 a_38516_n7844 0.285629f
C3175 a_33476_n20008 a_33564_n20052 0.285629f
C3176 a_29532_n20052 a_29980_n20052 0.012882f
C3177 a_34544_n2272 VDD 0.022627f
C3178 a_39724_n9509 a_40172_n9509 0.012222f
C3179 a_21772_n9860 a_21604_n10116 0.038564f
C3180 a_47812_n5896 VDD 0.211703f
C3181 a_26631_7 a_28352_n320 0.401636f
C3182 a_25831_n12996 VDD 0.715639f
C3183 a_21916_n1975 a_21828_n1931 0.495737f
C3184 a_45212_n15348 VDD 0.342281f
C3185 a_22164_n2760 a_24233_n3980 0.033345f
C3186 a_33452_n15781 a_33900_n15781 0.012882f
C3187 a_21692_2431 a_24628_1252 0.0215f
C3188 a_43196_n18484 VDD 0.316157f
C3189 a_47004_n16916 a_47116_n17349 0.026339f
C3190 a_26358_n4618 a_27190_n5112 0.106585f
C3191 a_24388_n4708 a_24180_n5112 0.027448f
C3192 a_21812_n6643 a_22052_n6980 0.068447f
C3193 a_39164_n18484 a_39276_n18917 0.026339f
C3194 a_23932_n18917 a_24380_n18917 0.013103f
C3195 a_42548_n7844 a_42996_n7844 0.013276f
C3196 a_43084_n9509 a_43444_n9412 0.087066f
C3197 a_27281_n16854 a_28435_n10599 0.211416f
C3198 a_43980_n6373 VDD 0.333977f
C3199 a_41740_n11077 a_42100_n10980 0.087066f
C3200 a_23564_n8292 a_23912_n15216 0.036226f
C3201 a_35120_n9412 VDD 0.013983f
C3202 a_23564_n11428 a_23360_n15233 0.05622f
C3203 a_35916_n12645 a_35828_n12548 0.285629f
C3204 a_44876_n12645 VDD 0.360805f
C3205 a_21772_n12996 a_22588_n16916 0.018617f
C3206 a_44316_n1236 a_44316_n1669 0.05841f
C3207 a_40172_n14213 a_40620_n14213 0.012001f
C3208 a_44428_n15781 VDD 0.321554f
C3209 a_35692_n15781 a_36052_n15684 0.087066f
C3210 a_46108_n2804 a_46220_n3237 0.026339f
C3211 a_42604_n2020 a_41684_n1976 0.014516f
C3212 a_25524_1243 a_26796_1515 0.05539f
C3213 a_35244_n18917 VDD 0.313885f
C3214 a_37036_n17349 a_36948_n17252 0.285629f
C3215 a_47116_n17349 a_47564_n17349 0.012882f
C3216 a_21692_n18917 a_21604_n18820 0.285629f
C3217 a_43892_n6276 a_44340_n6276 0.013276f
C3218 a_29612_n8292 a_30228_n8203 0.02278f
C3219 a_43196_n20052 a_43644_n20052 0.012882f
C3220 a_34460_n20052 a_34460_n20485 0.05841f
C3221 a_22876_n8988 a_23816_n8544 0.056721f
C3222 a_42636_n3237 VDD 0.315913f
C3223 a_46132_n9412 a_46580_n9412 0.013276f
C3224 a_28335_n10644 a_28927_n10160 0.108253f
C3225 a_33815_1384 VDD 1.32927f
C3226 a_37620_n12548 a_38068_n12548 0.013276f
C3227 a_46668_n12645 a_47028_n12548 0.087066f
C3228 a_21692_2431 a_28456_n364 0.014856f
C3229 a_21604_n13252 VDD 1.79896f
C3230 a_42636_n14213 a_42996_n14116 0.087066f
C3231 a_21604_n16872 VDD 0.221763f
C3232 a_46668_n15781 a_46580_n15684 0.285629f
C3233 a_25237_n4327 a_25423_n4328 0.356993f
C3234 a_37844_n15684 a_38292_n15684 0.013276f
C3235 a_33467_1116 a_34576_1204 0.019043f
C3236 a_30004_n18820 VDD 0.209535f
C3237 a_47564_n17349 a_47924_n17252 0.087066f
C3238 a_42636_n4805 a_42996_n4708 0.087066f
C3239 a_32332_n18917 a_32692_n18820 0.086635f
C3240 a_45772_n18917 a_46220_n18917 0.012882f
C3241 a_32543_n9032 a_32767_n9010 0.538085f
C3242 a_25860_n9032 a_25831_n11428 0.438126f
C3243 a_26271_n4306 VDD 0.314277f
C3244 a_38716_n7508 VDD 0.322794f
C3245 a_25627_n452 a_26736_n364 0.019043f
C3246 a_44004_n10600 VDD 0.2108f
C3247 a_28300_n15348 a_28212_n15303 0.104875f
C3248 a_44788_n14116 a_45236_n14116 0.013276f
C3249 a_35804_n16916 VDD 0.315469f
C3250 a_34860_n3189 a_33120_n3884 0.011422f
C3251 a_44340_n3140 a_44788_n3140 0.013276f
C3252 a_28836_376 a_28132_376 0.223572f
C3253 a_23396_n20008 VDD 0.207289f
C3254 a_23479_n5156 a_21812_n6643 0.017153f
C3255 a_22444_n5156 a_25612_n6679 0.079814f
C3256 a_22544_n4690 a_23949_n6724 0.075428f
C3257 a_31572_n17252 a_31684_n18440 0.026657f
C3258 a_39500_n6373 CLK 0.021787f
C3259 a_43532_n18917 a_43444_n18820 0.285629f
C3260 a_33497_n9032 a_34176_n6976 0.090554f
C3261 a_31656_n704 VDD 1.33837f
C3262 a_39164_n20485 a_39612_n20485 0.013103f
C3263 a_33868_n4240 VDD 0.298894f
C3264 a_30676_n7844 VDD 0.484919f
C3265 a_36164_n12168 a_35804_n12212 0.086905f
C3266 a_27167_n10808 VDD 0.566237f
C3267 a_47812_n13736 VDD 0.211703f
C3268 a_39636_n14116 a_39524_n15304 0.026657f
C3269 a_25160_n14816 a_25472_n14816 0.119687f
C3270 a_21692_2431 a_28671_n1976 0.492463f
C3271 a_46556_n16916 VDD 0.31705f
C3272 a_31684_n16872 a_32132_n16872 0.013276f
C3273 a_29532_n20052 VDD 0.333745f
C3274 a_38740_n17252 a_38628_n18440 0.026657f
C3275 a_32856_n7376 a_33308_n7376 0.026665f
C3276 a_42660_n7464 a_42300_n7508 0.087066f
C3277 a_21916_n1975 VDD 0.90957f
C3278 a_39612_n20485 a_39524_n20388 0.285629f
C3279 a_42748_n9076 a_43196_n9076 0.012882f
C3280 a_27281_n16854 a_28009_n12168 0.023696f
C3281 a_40420_n10600 a_40060_n10644 0.087066f
C3282 a_25573_n12167 a_25132_n16432 0.114867f
C3283 a_30781_n452 a_31405_n452 0.104193f
C3284 a_42548_n7844 VDD 0.205948f
C3285 a_42660_n12168 a_43108_n12168 0.013276f
C3286 a_38628_n12168 a_38716_n12212 0.285629f
C3287 a_42412_n101 a_42772_n4 0.086742f
C3288 a_32158_n12212 VDD 0.634898f
C3289 a_23564_n11428 a_25544_n16412 0.195196f
C3290 a_21772_n12996 a_21604_n15304 0.049878f
C3291 a_24233_n844 a_23816_n704 0.633318f
C3292 a_35604_n13736 a_35692_n13780 0.285629f
C3293 a_40172_n14213 VDD 0.315889f
C3294 a_33900_n15348 a_34348_n15348 0.013103f
C3295 a_46580_n14116 a_46468_n15304 0.026657f
C3296 a_47116_n17349 VDD 0.315469f
C3297 a_33015_n4284 a_33608_n4284 0.361958f
C3298 a_32359_n4372 a_33416_n4240 0.056721f
C3299 a_47028_n3140 a_46916_n4328 0.026657f
C3300 a_24631_n3588 a_28225_n4327 0.045855f
C3301 a_32579_769 a_32909_841 0.538085f
C3302 a_25975_n184 a_27032_51 0.056721f
C3303 a_43196_n20052 VDD 0.32959f
C3304 a_33028_n18440 a_33116_n18484 0.285629f
C3305 a_22220_n9860 a_23220_n7376 0.016849f
C3306 a_45684_n17252 a_45572_n18440 0.026657f
C3307 a_42212_n7464 CLK 0.043615f
C3308 a_47812_n7464 a_47900_n7508 0.285629f
C3309 a_46108_n7508 a_46556_n7508 0.012552f
C3310 a_34223_n1976 VDD 0.313315f
C3311 a_39524_n20388 a_39972_n20388 0.013276f
C3312 a_39748_2475 OUT[2] 0.023343f
C3313 a_34652_n11391 a_34350_n10980 0.391002f
C3314 a_46916_n10600 a_47364_n10600 0.013276f
C3315 a_45572_n10600 a_45660_n10644 0.285629f
C3316 a_32543_n9032 VDD 0.595077f
C3317 a_24464_n11680 VDD 0.040882f
C3318 a_31960_n13648 a_32412_n13648 0.026665f
C3319 a_27820_n16432 a_27192_n14286 0.712906f
C3320 a_40868_n13736 a_40956_n13780 0.285629f
C3321 a_29856_n1121 a_31968_n704 0.277491f
C3322 a_44788_n14116 VDD 0.22479f
C3323 a_41316_n15304 a_40956_n15348 0.087066f
C3324 a_47924_n17252 VDD 0.21239f
C3325 a_42660_n4328 a_42748_n4372 0.285629f
C3326 a_38716_n16916 a_39164_n16916 0.012882f
C3327 a_42660_n16872 a_42748_n16916 0.285629f
C3328 a_39164_n20485 VDD 0.302205f
C3329 a_46020_n5896 a_46108_n5940 0.285629f
C3330 a_47364_n5896 a_47812_n5896 0.013276f
C3331 a_26172_n20052 a_26620_n20052 0.012882f
C3332 a_40532_n18820 a_40420_n20008 0.026657f
C3333 a_22712_n7420 a_25831_n11428 0.067069f
C3334 a_47812_n1572 VDD 0.209236f
C3335 a_27281_n16854 a_22220_n12996 0.123445f
C3336 a_28624_n9394 a_28868_n9387 0.02407f
C3337 a_45212_n9076 a_45324_n9509 0.026339f
C3338 a_27281_n16854 a_27744_n12908 0.015095f
C3339 a_42748_n9076 VDD 0.315469f
C3340 a_24964_n14116 a_24516_n14475 0.209135f
C3341 a_21772_n12996 a_25132_n16432 0.015121f
C3342 a_22116_n12548 a_21892_n12952 0.013419f
C3343 a_42660_n12168 VDD 0.206217f
C3344 a_46468_n13736 a_46108_n13780 0.086905f
C3345 a_21772_n12996 a_22140_n15781 0.024807f
C3346 a_42884_n1192 a_42972_n1236 0.285629f
C3347 a_33900_n15348 VDD 0.296789f
C3348 a_46468_n15304 a_46556_n15348 0.285629f
C3349 a_27628_n3841 a_28583_n3140 0.02713f
C3350 a_40652_n1572 a_44316_n1669 0.015973f
C3351 a_36612_n18440 VDD 0.215061f
C3352 a_47812_n4328 a_47900_n4372 0.285629f
C3353 a_46108_n4372 a_46556_n4372 0.012552f
C3354 a_39524_n20388 VDD 0.207032f
C3355 a_42748_n18484 a_43196_n18484 0.012882f
C3356 a_45324_n7941 a_45772_n7941 0.012882f
C3357 a_33476_n20008 a_33116_n20052 0.087066f
C3358 a_38156_n7941 a_38516_n7844 0.087174f
C3359 a_47476_n18820 a_47364_n20008 0.026657f
C3360 a_47364_n5896 VDD 0.205948f
C3361 a_38380_n11077 a_38828_n11077 0.013103f
C3362 a_30871_n11728 a_30599_n12167 0.028982f
C3363 a_26736_n364 a_28352_n320 0.011851f
C3364 a_31235_n9860 VDD 0.331726f
C3365 a_29161_n14476 a_29056_n14432 0.116059f
C3366 a_44092_n13780 a_43980_n14213 0.026339f
C3367 a_47812_n15304 VDD 0.211703f
C3368 a_42748_n18484 VDD 0.315469f
C3369 a_36140_n17349 a_36588_n17349 0.012882f
C3370 a_43644_n4372 a_43532_n4805 0.026339f
C3371 a_30740_n7464 a_31936_n6592 0.09176f
C3372 a_43532_n6373 a_43980_n6373 0.012882f
C3373 a_30676_n7844 a_32543_n9032 0.055338f
C3374 a_39972_n20008 a_40420_n20008 0.013276f
C3375 a_25724_n14564 a_25412_n10600 0.04558f
C3376 a_43084_n9509 a_42996_n9412 0.285629f
C3377 a_43532_n6373 VDD 0.332233f
C3378 a_26239_n11428 a_26239_n12996 0.027963f
C3379 a_24684_n16432 a_25880_n11708 0.051043f
C3380 a_41740_n11077 a_41652_n10980 0.285629f
C3381 a_44428_n12645 a_44876_n12645 0.012882f
C3382 a_35468_n12645 a_35828_n12548 0.087174f
C3383 a_44428_n12645 VDD 0.321554f
C3384 a_21772_n12996 a_22140_n16916 0.032425f
C3385 a_43980_n15781 VDD 0.31896f
C3386 a_33588_n3461 a_36217_n3500 0.019043f
C3387 a_43980_n15781 a_44428_n15781 0.012882f
C3388 a_35692_n15781 a_35604_n15684 0.285629f
C3389 a_25524_1243 a_22096_376 0.10138f
C3390 a_34796_n18917 VDD 0.313885f
C3391 a_36588_n17349 a_36948_n17252 0.087066f
C3392 a_n199_2852 VIN 0.10575f
C3393 a_24492_n5156 a_25831_n11428 0.024618f
C3394 a_29612_n8292 a_28764_n8247 0.190361f
C3395 a_34796_n18917 a_35244_n18917 0.012882f
C3396 a_25972_n6276 a_33497_n9032 0.033758f
C3397 a_42188_n3237 VDD 0.315469f
C3398 a_25020_n11383 a_26239_n11428 0.236432f
C3399 a_33467_1116 VDD 0.475758f
C3400 a_28335_n10644 a_28437_n13705 0.043279f
C3401 a_26943_n7442 VDD 0.314737f
C3402 a_44340_n10980 a_44788_n10980 0.013276f
C3403 a_46668_n12645 a_46580_n12548 0.285629f
C3404 a_28121_n10980 a_29659_n14820 0.010009f
C3405 a_33812_n14116 a_34260_n14116 0.013276f
C3406 a_42636_n14213 a_42548_n14116 0.285629f
C3407 a_25237_n4327 a_23816_n3840 0.017205f
C3408 a_42188_n3237 a_42636_n3237 0.012882f
C3409 a_46220_n15781 a_46580_n15684 0.087066f
C3410 a_33467_1116 a_33815_1384 0.633318f
C3411 a_29556_n18820 VDD 0.20677f
C3412 a_47564_n17349 a_47476_n17252 0.285629f
C3413 a_36948_n17252 a_37396_n17252 0.013276f
C3414 a_42636_n4805 a_42548_n4708 0.285629f
C3415 a_25612_n6679 a_33308_n7376 0.01791f
C3416 a_32332_n18917 a_32244_n18820 0.285629f
C3417 a_26047_n4328 VDD 0.587353f
C3418 a_25724_n14564 a_24964_n14116 0.380796f
C3419 a_39636_n9412 a_39524_n10600 0.026657f
C3420 a_38268_n7508 VDD 0.357068f
C3421 a_38292_n10980 a_38180_n12168 0.026657f
C3422 a_24684_n16432 a_26239_n12996 0.323786f
C3423 a_24964_n14116 a_27639_n12537 0.041213f
C3424 a_25627_n452 a_25975_n184 0.633318f
C3425 a_43556_n10600 VDD 0.209225f
C3426 a_22600_n12124 a_22140_n15348 0.033245f
C3427 a_47452_n1669 a_47900_n1669 0.012001f
C3428 a_35356_n16916 VDD 0.315469f
C3429 a_34000_n3140 a_33120_n3884 0.014454f
C3430 a_34708_n15684 a_34820_n16872 0.026657f
C3431 a_22052_n4708 a_28144_n4708 0.026401f
C3432 a_31324_n4372 a_30104_n1148 0.017545f
C3433 a_41616_1564 a_42168_1564 0.361958f
C3434 a_41864_1394 a_41964_1564 0.11204f
C3435 a_22948_n20008 VDD 0.205626f
C3436 a_28836_376 a_28492_332 0.038295f
C3437 a_24492_n5156 a_23619_n6724 0.047355f
C3438 a_47028_n4708 a_47476_n4708 0.013276f
C3439 a_46580_n6276 a_46468_n7464 0.026657f
C3440 a_29556_n18820 a_30004_n18820 0.013276f
C3441 a_43084_n18917 a_43444_n18820 0.087066f
C3442 a_32073_n844 VDD 0.479301f
C3443 a_39972_n9032 a_40420_n9032 0.013276f
C3444 a_29532_n10311 a_32581_n9860 0.13538f
C3445 a_33672_n10112 a_33984_n10112 0.119687f
C3446 a_46580_n9412 a_46468_n10600 0.026657f
C3447 a_27281_n16854 a_28300_n15348 0.014131f
C3448 a_35816_n174 VDD 0.432917f
C3449 a_35716_n12168 a_35804_n12212 0.285629f
C3450 a_41204_n12548 a_41316_n13736 0.026657f
C3451 a_47364_n13736 VDD 0.205948f
C3452 a_27404_n14990 a_27852_n14990 0.237602f
C3453 a_25577_n14956 a_25472_n14816 0.116059f
C3454 a_22500_n1976 a_23954_n2020 0.015579f
C3455 a_46108_n16916 VDD 0.318654f
C3456 a_23816_n3840 a_24128_n3840 0.119687f
C3457 a_26047_n4328 a_26271_n4306 0.538085f
C3458 a_39860_n3140 a_39972_n4328 0.026657f
C3459 a_42100_n15684 a_42212_n16872 0.026657f
C3460 a_36612_n20008 VDD 0.215061f
C3461 a_24828_n18484 a_25276_n18484 0.012222f
C3462 a_38268_n7508 a_38716_n7508 0.012882f
C3463 a_26420_n18820 a_26532_n20008 0.026657f
C3464 a_42212_n7464 a_42300_n7508 0.285629f
C3465 a_47900_n1236 VDD 0.318055f
C3466 a_39164_n20485 a_39524_n20388 0.087174f
C3467 a_43556_n10600 a_44004_n10600 0.013276f
C3468 a_23564_n8292 a_24128_n13248 0.03746f
C3469 a_39972_n10600 a_40060_n10644 0.285629f
C3470 a_25573_n12167 a_25559_n12548 0.032381f
C3471 a_24628_n363 VDD 0.521221f
C3472 a_42100_n7844 VDD 0.205948f
C3473 a_26431_n12168 a_26983_n12728 0.021389f
C3474 a_38628_n12168 a_38268_n12212 0.087066f
C3475 a_24964_n14116 a_25237_n13735 0.025279f
C3476 a_35604_n13736 a_35244_n13780 0.086905f
C3477 a_39724_n14213 VDD 0.319134f
C3478 a_23004_n2332 a_22772_n1104 0.024225f
C3479 a_46668_n17349 VDD 0.318039f
C3480 a_22052_n4708 a_27190_n5112 0.010516f
C3481 a_35356_n16916 a_35804_n16916 0.012222f
C3482 a_33120_n3884 a_33608_n4284 0.08126f
C3483 a_42748_n20052 VDD 0.328902f
C3484 a_42772_n5896 a_43220_n5896 0.013276f
C3485 a_22220_n9860 a_24576_n6976 0.051132f
C3486 a_33028_n18440 a_32668_n18484 0.087066f
C3487 a_41764_n7464 CLK 0.013118f
C3488 a_33364_n18820 a_33476_n20008 0.026657f
C3489 a_22948_n20008 a_23396_n20008 0.013276f
C3490 a_47812_n7464 a_47452_n7508 0.086635f
C3491 a_33999_n1400 VDD 0.578623f
C3492 a_22264_n10556 a_23949_n9860 0.013823f
C3493 a_23619_n9860 a_24965_n9860 0.042679f
C3494 a_48012_n4805 VDD 0.343411f
C3495 a_45572_n10600 a_45212_n10644 0.086905f
C3496 a_34652_n11391 a_35064_n11383 0.018413f
C3497 a_31919_n9032 VDD 0.7306f
C3498 a_28121_n10980 a_29479_n13735 0.045959f
C3499 a_44540_n12212 a_45124_n12168 0.016748f
C3500 a_40868_n13736 a_40508_n13780 0.087066f
C3501 a_32073_n844 a_31656_n704 0.633318f
C3502 a_44340_n14116 VDD 0.212126f
C3503 a_40868_n15304 a_40956_n15348 0.285629f
C3504 a_28736_1944 a_22164_n2760 0.027646f
C3505 a_31324_n4372 a_22820_n2804 0.023741f
C3506 a_47476_n17252 VDD 0.206217f
C3507 a_30428_n16916 a_30316_n17349 0.026339f
C3508 a_42660_n16872 a_42300_n16916 0.087066f
C3509 a_42660_n4328 a_42300_n4372 0.086905f
C3510 a_38716_n20485 VDD 0.304516f
C3511 a_24380_n18484 a_24380_n18917 0.05841f
C3512 a_39524_n18440 a_39972_n18440 0.013276f
C3513 a_46020_n5896 a_45660_n5940 0.086905f
C3514 a_45660_n7508 a_45772_n7941 0.026339f
C3515 a_47364_n1572 VDD 0.203482f
C3516 a_42748_n10644 a_42636_n11077 0.026339f
C3517 a_27281_n16854 a_26983_n12728 0.051991f
C3518 a_42300_n9076 VDD 0.315469f
C3519 a_21872_n12530 a_21892_n12952 0.576301f
C3520 a_39164_n12212 a_39052_n12645 0.026339f
C3521 a_42212_n12168 VDD 0.206217f
C3522 a_47364_n13736 a_47812_n13736 0.013276f
C3523 a_46020_n13736 a_46108_n13780 0.285629f
C3524 a_21772_n12996 a_21692_n15781 0.057791f
C3525 a_33452_n15348 VDD 0.296789f
C3526 a_46468_n15304 a_46108_n15348 0.086905f
C3527 a_41180_n2804 a_41628_n2804 0.013103f
C3528 a_40652_n1572 a_43868_n1669 0.014145f
C3529 a_36164_n18440 VDD 0.206217f
C3530 a_47812_n4328 a_47452_n4372 0.086635f
C3531 a_47812_n16872 a_47900_n16916 0.285629f
C3532 a_37372_n16916 a_37484_n17349 0.026339f
C3533 a_46108_n16916 a_46556_n16916 0.012552f
C3534 a_44452_376 a_44540_332 0.285629f
C3535 a_39076_n20388 VDD 0.208947f
C3536 a_31772_n18484 a_31884_n18917 0.026339f
C3537 a_33028_n20008 a_33116_n20052 0.285629f
C3538 a_38156_n7941 a_38068_n7844 0.285629f
C3539 a_29732_n2760 VDD 0.014136f
C3540 a_39276_n9509 a_39724_n9509 0.013103f
C3541 a_46916_n5896 VDD 0.205962f
C3542 a_26631_7 a_28456_n364 0.340745f
C3543 a_27224_n62 a_27484_n4 0.66083f
C3544 a_42636_n17349 CLK 0.01698f
C3545 a_30472_n9815 VDD 0.457758f
C3546 a_28744_n14432 a_29056_n14432 0.119687f
C3547 a_47364_n15304 VDD 0.205948f
C3548 a_39357_n2228 a_39500_n3237 0.031039f
C3549 a_42300_n18484 VDD 0.315469f
C3550 a_46556_n16916 a_46668_n17349 0.026339f
C3551 a_38716_n18484 a_38828_n18917 0.026339f
C3552 a_23484_n18917 a_23932_n18917 0.013103f
C3553 a_31341_n8292 a_30900_n9032 0.03774f
C3554 a_42100_n7844 a_42548_n7844 0.013276f
C3555 a_30676_n7844 a_31919_n9032 0.463602f
C3556 a_42636_n9509 a_42996_n9412 0.087066f
C3557 a_25084_1564 VDD 1.77402f
C3558 a_43084_n6373 VDD 0.328902f
C3559 a_41292_n11077 a_41652_n10980 0.087066f
C3560 a_23564_n8292 a_24220_n15260 0.02323f
C3561 a_28335_n10644 VDD 0.404293f
C3562 a_22264_n13692 a_22364_n13648 0.09301f
C3563 a_35468_n12645 a_35380_n12548 0.285629f
C3564 a_43980_n12645 VDD 0.31896f
C3565 a_28671_n1976 a_29295_n1400 0.104193f
C3566 a_21772_n12996 a_21692_n16916 0.030287f
C3567 a_39724_n14213 a_40172_n14213 0.012882f
C3568 a_43532_n15781 VDD 0.317216f
C3569 a_45660_n2804 a_45772_n3237 0.026339f
C3570 a_33588_n3461 a_35800_n3456 0.042802f
C3571 a_35244_n15781 a_35604_n15684 0.087066f
C3572 a_25524_1243 a_25936_1564 0.536965f
C3573 a_24628_1252 a_22096_376 0.011013f
C3574 a_25084_1564 a_33815_1384 0.023168f
C3575 a_34348_n18917 VDD 0.313885f
C3576 a_36588_n17349 a_36500_n17252 0.285629f
C3577 a_46668_n17349 a_47116_n17349 0.012882f
C3578 a_47900_n18484 a_48012_n18917 0.026339f
C3579 a_43444_n6276 a_43892_n6276 0.013276f
C3580 a_22016_n8961 a_23816_n8544 0.510371f
C3581 a_34012_n20052 a_34012_n20485 0.05841f
C3582 a_42748_n20052 a_43196_n20052 0.012882f
C3583 a_25972_n6276 a_33672_n10112 0.011277f
C3584 a_41740_n3237 VDD 0.315669f
C3585 a_45684_n9412 a_46132_n9412 0.013276f
C3586 a_27484_n4 VDD 0.298894f
C3587 a_26719_n7464 VDD 0.578598f
C3588 a_26239_n11428 VDD 0.501748f
C3589 a_30340_n12548 a_30555_n13780 0.02132f
C3590 a_37172_n12548 a_37620_n12548 0.013276f
C3591 a_46220_n12645 a_46580_n12548 0.087066f
C3592 a_47924_n12548 VDD 0.21239f
C3593 a_42188_n14213 a_42548_n14116 0.087066f
C3594 a_33999_n1400 a_34223_n1976 0.538085f
C3595 a_47924_n15684 VDD 0.21239f
C3596 a_46220_n15781 a_46132_n15684 0.285629f
C3597 a_25237_n4327 a_24233_n3980 0.111804f
C3598 a_37396_n15684 a_37844_n15684 0.013276f
C3599 a_29108_n18820 VDD 0.209318f
C3600 a_25237_n5895 a_25412_n5895 0.134967f
C3601 a_42188_n4805 a_42548_n4708 0.087066f
C3602 a_47116_n17349 a_47476_n17252 0.087066f
C3603 a_24631_n3588 a_25972_n6276 0.010975f
C3604 a_45324_n18917 a_45772_n18917 0.012882f
C3605 a_21812_n6643 a_24752_n8292 0.015037f
C3606 a_31884_n18917 a_32244_n18820 0.087066f
C3607 a_25573_n12167 a_28225_n9031 0.188851f
C3608 a_31919_n9032 a_32543_n9032 0.104193f
C3609 a_25423_n4328 VDD 0.707955f
C3610 a_23524_464 VDD 0.01368f
C3611 a_37820_n7508 VDD 0.324073f
C3612 a_24684_n16432 a_25831_n12996 0.110961f
C3613 a_24964_n14116 a_25132_n16432 0.195831f
C3614 a_26547_n12951 a_25559_n12548 0.104402f
C3615 a_43108_n10600 VDD 0.206217f
C3616 a_36500_n13736 VDD 0.216152f
C3617 a_44340_n14116 a_44788_n14116 0.013276f
C3618 a_34908_n16916 VDD 0.315469f
C3619 a_43892_n3140 a_44340_n3140 0.013276f
C3620 a_30555_n2729 a_32132_n4708 0.13071f
C3621 a_27988_n20388 a_27988_n17252 0.011945f
C3622 a_42604_n2020 a_42436_n2760 0.036074f
C3623 a_41616_1564 a_41964_1564 0.401636f
C3624 a_22500_n20008 VDD 0.203482f
C3625 a_47476_n17252 a_47924_n17252 0.013276f
C3626 a_23887_n5156 a_23619_n6724 0.054704f
C3627 a_31124_n17252 a_31236_n18440 0.026657f
C3628 a_43084_n18917 a_42996_n18820 0.285629f
C3629 a_24492_n5156 a_29992_n11150 0.012846f
C3630 a_29532_n10311 a_32189_n9860 0.070487f
C3631 a_26844_n20485 a_26756_n20388 0.285629f
C3632 a_38716_n20485 a_39164_n20485 0.013103f
C3633 a_34736_n3840 VDD 0.010384f
C3634 a_32424_n10512 a_32628_n10512 0.66083f
C3635 a_34089_n10252 a_33984_n10112 0.116059f
C3636 a_25020_n11383 a_25559_n10980 0.013683f
C3637 a_35716_n12168 a_35356_n12212 0.086905f
C3638 a_24684_n16432 VDD 0.771812f
C3639 a_46916_n13736 VDD 0.205962f
C3640 a_47364_n1572 a_47812_n1572 0.013276f
C3641 a_39188_n14116 a_39076_n15304 0.026657f
C3642 a_22500_n1976 a_23542_n1754 0.086212f
C3643 a_45660_n16916 VDD 0.320877f
C3644 a_31236_n16872 a_31684_n16872 0.013276f
C3645 a_24233_n3980 a_24128_n3840 0.116059f
C3646 a_36164_n20008 VDD 0.206217f
C3647 a_24041_816 a_24913_864 0.152869f
C3648 a_38292_n17252 a_38180_n18440 0.026657f
C3649 a_30036_n7464 a_30228_n8203 0.011489f
C3650 a_42212_n7464 a_41852_n7508 0.087066f
C3651 a_30396_n7508 a_31011_n8292 0.214895f
C3652 a_40084_n18820 a_40532_n18820 0.013276f
C3653 a_21812_n6643 a_21872_n9394 0.040152f
C3654 a_47452_n1236 VDD 0.296789f
C3655 a_42300_n9076 a_42748_n9076 0.012882f
C3656 a_25860_n9032 a_25724_n14564 0.033439f
C3657 a_39164_n20485 a_39076_n20388 0.285629f
C3658 a_22220_n9860 VDD 1.49722f
C3659 a_39972_n10600 a_39612_n10644 0.087066f
C3660 a_41652_n7844 VDD 0.205948f
C3661 a_42212_n12168 a_42660_n12168 0.013276f
C3662 a_46132_n4 VDD 0.2106f
C3663 a_26563_n12212 a_26983_n12728 0.029196f
C3664 a_24964_n14116 a_23816_n13248 0.019083f
C3665 a_38180_n12168 a_38268_n12212 0.285629f
C3666 a_47924_n12548 a_47812_n13736 0.026657f
C3667 a_35156_n13736 a_35244_n13780 0.285629f
C3668 a_22016_n1121 a_24128_n704 0.277491f
C3669 a_24631_n3588 a_31405_n452 0.038105f
C3670 a_39276_n14213 VDD 0.320782f
C3671 a_46132_n14116 a_46020_n15304 0.026657f
C3672 a_33452_n15348 a_33900_n15348 0.013103f
C3673 a_27452_n2716 a_27348_n2672 0.11011f
C3674 a_46220_n17349 VDD 0.31977f
C3675 a_33120_n3884 a_33015_n4284 0.536965f
C3676 a_46580_n3140 a_46468_n4328 0.026657f
C3677 a_32359_n4372 a_32911_n4240 0.119687f
C3678 a_42300_n20052 VDD 0.328902f
C3679 a_45236_n17252 a_45124_n18440 0.026657f
C3680 a_36164_n18440 a_36612_n18440 0.013276f
C3681 a_32580_n18440 a_32668_n18484 0.285629f
C3682 a_22444_n5156 a_33048_n7420 0.01252f
C3683 a_41316_n7464 CLK 0.012286f
C3684 a_45660_n7508 a_46108_n7508 0.012552f
C3685 a_47364_n7464 a_47452_n7508 0.285629f
C3686 a_39076_n20388 a_39524_n20388 0.013276f
C3687 a_21772_n9860 a_24965_n9860 0.01999f
C3688 a_23479_n5156 a_26470_n13736 0.05472f
C3689 a_29532_n10311 a_30808_n10116 0.010901f
C3690 a_47564_n4805 VDD 0.315469f
C3691 a_45124_n10600 a_45212_n10644 0.285629f
C3692 a_46468_n10600 a_46916_n10600 0.013276f
C3693 a_30900_n9032 VDD 0.615023f
C3694 a_27279_n12146 VDD 0.316607f
C3695 a_40420_n13736 a_40508_n13780 0.285629f
C3696 a_44004_n13736 a_44452_n13736 0.013276f
C3697 a_43892_n14116 VDD 0.210071f
C3698 a_40868_n15304 a_40508_n15348 0.087066f
C3699 a_34248_n3310 a_33588_n3461 0.09725f
C3700 a_22500_n1976 a_22164_n2760 0.408954f
C3701 a_30104_n1148 a_30204_n1104 0.088f
C3702 a_47028_n17252 VDD 0.206217f
C3703 a_42212_n16872 a_42300_n16916 0.285629f
C3704 a_42212_n4328 a_42300_n4372 0.285629f
C3705 a_38268_n16916 a_38716_n16916 0.012882f
C3706 a_38268_n20485 VDD 0.336417f
C3707 a_46916_n5896 a_47364_n5896 0.013276f
C3708 a_45572_n5896 a_45660_n5940 0.285629f
C3709 a_25724_n20052 a_26172_n20052 0.012882f
C3710 a_40084_n18820 a_39972_n20008 0.026657f
C3711 a_46916_n1572 VDD 0.203495f
C3712 a_42748_n13780 CLK 0.012909f
C3713 a_22220_n12996 a_21872_n12530 0.428867f
C3714 a_41852_n9076 VDD 0.315469f
C3715 a_28300_n15348 a_34708_n13736 0.024586f
C3716 a_137_4292 VDD 0.542539f
C3717 a_41764_n12168 VDD 0.206217f
C3718 a_46020_n13736 a_45660_n13780 0.086905f
C3719 a_36588_n13780 a_36588_n14213 0.05841f
C3720 a_22600_n12124 a_23484_n16916 0.011887f
C3721 a_33004_n15348 VDD 0.331004f
C3722 a_46020_n15304 a_46108_n15348 0.285629f
C3723 a_32020_n2276 a_33588_n3461 0.138296f
C3724 a_47364_n15304 a_47812_n15304 0.013276f
C3725 a_40652_n1572 a_43420_n1669 0.013445f
C3726 a_35716_n18440 VDD 0.206217f
C3727 a_47364_n4328 a_47452_n4372 0.285629f
C3728 a_47812_n16872 a_47452_n16916 0.086635f
C3729 a_45660_n4372 a_46108_n4372 0.012552f
C3730 a_38628_n20388 VDD 0.211896f
C3731 a_42300_n18484 a_42748_n18484 0.012882f
C3732 a_47028_n18820 a_46916_n20008 0.026657f
C3733 a_37708_n7941 a_38068_n7844 0.087174f
C3734 a_33028_n20008 a_32668_n20052 0.087066f
C3735 a_44876_n7941 a_45324_n7941 0.012882f
C3736 a_46468_n5896 VDD 0.209055f
C3737 a_37932_n11077 a_38380_n11077 0.013103f
C3738 a_30871_n11728 a_31760_n12168 0.015767f
C3739 a_26736_n364 a_28456_n364 0.107654f
C3740 a_42188_n17349 CLK 0.047331f
C3741 a_28624_n9394 VDD 0.483158f
C3742 a_24573_n12996 VDD 0.8506f
C3743 a_43644_n13780 a_43532_n14213 0.026339f
C3744 a_26944_n14116 a_28752_n15348 0.032605f
C3745 a_28744_n14432 a_29161_n14476 0.633318f
C3746 a_46916_n15304 VDD 0.205962f
C3747 a_22164_n2760 a_22568_n4240 0.025463f
C3748 a_41852_n18484 VDD 0.315469f
C3749 a_35692_n17349 a_36140_n17349 0.012882f
C3750 a_43196_n4372 a_43084_n4805 0.026339f
C3751 a_43084_n6373 a_43532_n6373 0.012882f
C3752 a_39524_n20008 a_39972_n20008 0.013276f
C3753 a_22712_n7420 a_25724_n14564 0.01129f
C3754 a_30676_n7844 a_30900_n9032 0.024712f
C3755 a_27281_n16854 a_28927_n10160 0.022614f
C3756 a_42636_n9509 a_42548_n9412 0.285629f
C3757 a_22220_n12996 a_27485_n10068 0.02834f
C3758 a_42636_n6373 VDD 0.328902f
C3759 a_41292_n11077 a_41204_n10980 0.285629f
C3760 a_23564_n8292 a_23608_n15260 0.061791f
C3761 a_35020_n12645 a_35380_n12548 0.087174f
C3762 a_43980_n12645 a_44428_n12645 0.012882f
C3763 a_43532_n12645 VDD 0.317216f
C3764 a_43556_n661 a_43868_n1669 0.029777f
C3765 a_43084_n15781 VDD 0.313885f
C3766 a_35244_n15781 a_35156_n15684 0.285629f
C3767 a_43532_n15781 a_43980_n15781 0.012882f
C3768 a_33900_n18917 VDD 0.313885f
C3769 a_36140_n17349 a_36500_n17252 0.087066f
C3770 a_23479_n5156 a_25831_n11428 0.051077f
C3771 a_34348_n18917 a_34796_n18917 0.012882f
C3772 a_22364_n8944 a_22568_n8944 0.048436f
C3773 a_22016_n8961 a_24233_n8684 0.020455f
C3774 a_21604_n8548 a_23816_n8544 0.042802f
C3775 a_29532_n10311 a_25831_n11428 0.031933f
C3776 a_41292_n3237 VDD 0.321686f
C3777 a_31856_1248 VDD 0.025398f
C3778 a_26095_n7464 VDD 0.713535f
C3779 a_43892_n10980 a_44340_n10980 0.013276f
C3780 a_25500_n10644 VDD 0.3278f
C3781 a_46220_n12645 a_46132_n12548 0.285629f
C3782 a_47476_n12548 VDD 0.206217f
C3783 a_33364_n14116 a_33812_n14116 0.013276f
C3784 a_42188_n14213 a_42100_n14116 0.285629f
C3785 a_47476_n15684 VDD 0.206217f
C3786 a_41740_n3237 a_42188_n3237 0.012882f
C3787 a_45772_n15781 a_46132_n15684 0.087066f
C3788 a_28660_n18820 VDD 0.206648f
C3789 a_44004_n1192 a_40652_n1572 0.033614f
C3790 a_36500_n17252 a_36948_n17252 0.013276f
C3791 a_42188_n4805 a_42100_n4708 0.285629f
C3792 a_47116_n17349 a_47028_n17252 0.285629f
C3793 a_24672_n11339 a_25412_n5895 0.132424f
C3794 a_48012_n101 VDD 0.32473f
C3795 a_31884_n18917 a_31796_n18820 0.285629f
C3796 a_21812_n6643 a_23564_n8292 0.017826f
C3797 a_39412_n6276 a_39524_n7464 0.026657f
C3798 a_26719_n7464 a_26943_n7442 0.538085f
C3799 a_26396_n20485 a_26844_n20485 0.012552f
C3800 a_23816_n3840 VDD 1.37609f
C3801 a_27281_n16854 a_29332_n11301 0.010905f
C3802 a_39188_n9412 a_39076_n10600 0.026657f
C3803 a_23728_464 VDD 0.271996f
C3804 a_42748_n15348 CLK 0.012909f
C3805 a_37372_n7508 VDD 0.329356f
C3806 a_24964_n14116 a_25559_n12548 0.096413f
C3807 a_37844_n10980 a_37732_n12168 0.026657f
C3808 a_26431_n12168 a_25880_n11708 0.228163f
C3809 a_42660_n10600 VDD 0.206217f
C3810 a_36052_n13736 VDD 0.208855f
C3811 a_41292_n1669 a_41204_n1572 0.285629f
C3812 a_47004_n1669 a_47452_n1669 0.012222f
C3813 a_34460_n16916 VDD 0.315469f
C3814 a_34260_n15684 a_34372_n16872 0.026657f
C3815 a_41616_1564 a_42476_1515 0.882105f
C3816 a_22052_n20008 VDD 0.203482f
C3817 a_46580_n4708 a_47028_n4708 0.013276f
C3818 a_46132_n6276 a_46020_n7464 0.026657f
C3819 a_24492_n5156 a_25724_n14564 0.031976f
C3820 a_29108_n18820 a_29556_n18820 0.013276f
C3821 a_42636_n18917 a_42996_n18820 0.087066f
C3822 VDD OUT[0] 0.932626f
C3823 a_26396_n20485 a_26756_n20388 0.086905f
C3824 a_39524_n9032 a_39972_n9032 0.013276f
C3825 a_46132_n9412 a_46020_n10600 0.026657f
C3826 a_29176_n7819 VDD 0.021926f
C3827 a_35268_n12168 a_35356_n12212 0.285629f
C3828 a_25559_n10980 VDD 0.971207f
C3829 a_46468_n13736 VDD 0.209055f
C3830 a_23912_n15216 a_24116_n15216 0.66083f
C3831 a_22500_n1976 a_22918_n2020 0.056951f
C3832 a_45212_n16916 VDD 0.342281f
C3833 a_41652_n15684 a_41764_n16872 0.026657f
C3834 a_25423_n4328 a_26047_n4328 0.104193f
C3835 a_39412_n3140 a_39524_n4328 0.026657f
C3836 a_23136_447 a_25137_864 0.056679f
C3837 a_35716_n20008 VDD 0.206217f
C3838 a_28436_n18440 a_28524_n18484 0.285629f
C3839 a_24380_n18484 a_24828_n18484 0.013103f
C3840 a_25972_n18820 a_26084_n20008 0.026657f
C3841 a_33048_n7420 a_33308_n7376 0.66083f
C3842 a_37820_n7508 a_38268_n7508 0.012882f
C3843 a_41764_n7464 a_41852_n7508 0.285629f
C3844 a_47004_n1236 VDD 0.296789f
C3845 a_38716_n20485 a_39076_n20388 0.087174f
C3846 a_26308_n20388 a_26756_n20388 0.013276f
C3847 a_30900_n9032 a_31235_n9860 0.028277f
C3848 a_39524_n10600 a_39612_n10644 0.285629f
C3849 a_43108_n10600 a_43556_n10600 0.013276f
C3850 a_30451_n452 a_30781_n452 0.538085f
C3851 a_41204_n7844 VDD 0.227793f
C3852 a_26563_n12212 a_26635_n12996 0.027826f
C3853 a_38180_n12168 a_37820_n12212 0.087066f
C3854 a_24964_n14116 a_24233_n13388 0.041136f
C3855 a_48012_n11077 VDD 0.343411f
C3856 a_22600_n12124 a_23036_n15781 0.016383f
C3857 a_35156_n13736 a_34796_n13780 0.086905f
C3858 a_24631_n3588 a_30781_n452 0.067764f
C3859 a_38828_n14213 VDD 0.323023f
C3860 a_36500_n15304 a_36588_n15348 0.285629f
C3861 a_45772_n17349 VDD 0.321879f
C3862 a_34908_n16916 a_35356_n16916 0.012552f
C3863 a_31787_n3969 a_32911_n4240 0.116229f
C3864 a_41852_n20052 VDD 0.328902f
C3865 a_42324_n5896 a_42772_n5896 0.013276f
C3866 a_22444_n5156 a_32455_n7420 0.017956f
C3867 a_32580_n18440 a_32220_n18484 0.087066f
C3868 a_40868_n7464 CLK 0.010636f
C3869 a_47364_n7464 a_47004_n7508 0.086742f
C3870 a_22500_n20008 a_22948_n20008 0.013276f
C3871 a_23479_n5156 a_26266_n13736 0.010853f
C3872 a_23619_n9860 a_23949_n9860 0.538085f
C3873 a_36388_1944 OUT[2] 0.051004f
C3874 a_47116_n4805 VDD 0.315469f
C3875 a_31760_n12168 a_32413_n12996 0.017571f
C3876 a_44092_n12212 a_44540_n12212 0.012001f
C3877 a_27055_n12168 VDD 0.580765f
C3878 a_32152_n13692 a_32412_n13648 0.66083f
C3879 a_40420_n13736 a_40060_n13780 0.087066f
C3880 a_43444_n14116 VDD 0.208665f
C3881 a_34232_n2272 a_34544_n2272 0.119687f
C3882 a_40420_n15304 a_40508_n15348 0.285629f
C3883 a_27852_n14990 a_27709_n16132 0.023521f
C3884 a_44004_n15304 a_44452_n15304 0.013276f
C3885 a_28736_1944 a_22820_n2804 0.033416f
C3886 a_46580_n17252 VDD 0.209016f
C3887 a_42212_n4328 a_41852_n4372 0.087174f
C3888 a_42212_n16872 a_41852_n16916 0.087066f
C3889 a_37820_n20485 VDD 0.30591f
C3890 a_23932_n18484 a_23932_n18917 0.05841f
C3891 a_39076_n18440 a_39524_n18440 0.013276f
C3892 a_45572_n5896 a_45212_n5940 0.086905f
C3893 a_45212_n7508 a_45324_n7941 0.026339f
C3894 a_46468_n1572 VDD 0.206589f
C3895 a_42300_n13780 CLK 0.048577f
C3896 a_42300_n10644 a_42188_n11077 0.026339f
C3897 a_41404_n9076 VDD 0.315469f
C3898 a_38716_n12212 a_38604_n12645 0.026339f
C3899 a_23564_n11428 a_24516_n14475 0.013935f
C3900 a_21772_n12996 a_21892_n12952 0.392261f
C3901 a_28300_n15348 a_29479_n13735 0.013979f
C3902 a_41316_n12168 VDD 0.206217f
C3903 a_46916_n13736 a_47364_n13736 0.013276f
C3904 a_26431_n1192 a_26271_n1400 0.018117f
C3905 a_45572_n13736 a_45660_n13780 0.285629f
C3906 a_22600_n12124 a_23036_n16916 0.012134f
C3907 a_28212_n15303 VDD 0.629541f
C3908 a_46020_n15304 a_45660_n15348 0.086905f
C3909 a_40732_n2804 a_41180_n2804 0.013103f
C3910 a_27628_n3841 a_25600_n5895 0.04998f
C3911 a_22164_n2760 a_22052_n4708 0.013689f
C3912 a_40652_n1572 a_42244_n1572 0.037788f
C3913 a_35268_n18440 VDD 0.206217f
C3914 a_47364_n4328 a_47004_n4372 0.086742f
C3915 a_47364_n16872 a_47452_n16916 0.285629f
C3916 a_45660_n16916 a_46108_n16916 0.012552f
C3917 a_38180_n20388 VDD 0.243302f
C3918 a_31324_n18484 a_31436_n18917 0.026339f
C3919 a_25524_n6635 a_25972_n6276 0.195905f
C3920 a_36164_n20008 a_36612_n20008 0.013276f
C3921 a_32580_n20008 a_32668_n20052 0.285629f
C3922 a_37708_n7941 a_37620_n7844 0.285629f
C3923 a_34232_n2272 VDD 1.31068f
C3924 a_23479_n5156 a_26532_n14437 0.06446f
C3925 a_27281_n16854 a_25020_n11383 0.525949f
C3926 a_38828_n9509 a_39276_n9509 0.013103f
C3927 a_46020_n5896 VDD 0.210736f
C3928 a_29800_n9815 VDD 0.440108f
C3929 a_47900_n12212 a_48012_n12645 0.026339f
C3930 a_31789_n12996 a_32413_n12996 0.104193f
C3931 a_23949_n12996 VDD 0.569823f
C3932 a_47452_n1236 a_47900_n1236 0.012001f
C3933 a_46468_n15304 VDD 0.209055f
C3934 a_41404_n18484 VDD 0.315469f
C3935 a_46108_n16916 a_46220_n17349 0.026339f
C3936 a_22220_n9860 a_24836_n4708 0.012522f
C3937 a_22968_n6679 a_22052_n6980 0.014976f
C3938 a_23036_n18917 a_23484_n18917 0.013103f
C3939 a_38268_n18484 a_38380_n18917 0.026339f
C3940 a_41652_n7844 a_42100_n7844 0.013276f
C3941 a_47900_n2804 VDD 0.335152f
C3942 a_31324_n4372 VDD 1.45034f
C3943 a_22220_n12996 a_26861_n10135 0.011824f
C3944 a_27281_n16854 a_28437_n13705 0.029299f
C3945 a_42188_n9509 a_42548_n9412 0.087066f
C3946 a_42188_n6373 VDD 0.328902f
C3947 a_27167_n10808 a_27055_n12168 0.026651f
C3948 a_23564_n8292 a_23360_n15233 0.037754f
C3949 a_40620_n11077 a_41204_n10980 0.016748f
C3950 a_42548_n17252 CLK 0.029747f
C3951 a_35020_n12645 a_34932_n12548 0.285629f
C3952 a_22264_n13692 a_22016_n13665 0.348136f
C3953 a_43084_n12645 VDD 0.313885f
C3954 a_39276_n14213 a_39724_n14213 0.012882f
C3955 a_42636_n15781 VDD 0.313885f
C3956 a_33588_n3461 a_34552_n3140 0.08126f
C3957 a_45212_n2804 a_45324_n3237 0.026339f
C3958 a_34796_n15781 a_35156_n15684 0.087066f
C3959 a_33452_n18917 VDD 0.318502f
C3960 a_36140_n17349 a_36052_n17252 0.285629f
C3961 a_46220_n17349 a_46668_n17349 0.012882f
C3962 a_42996_n6276 a_43444_n6276 0.013276f
C3963 a_47452_n18484 a_47564_n18917 0.026339f
C3964 a_30740_n7464 a_30036_n7464 0.22378f
C3965 a_29532_n10311 a_34092_n9076 0.696952f
C3966 a_33564_n20052 a_33564_n20485 0.05841f
C3967 a_42300_n20052 a_42748_n20052 0.012882f
C3968 a_21604_n8548 a_24233_n8684 0.019043f
C3969 a_22876_n8988 a_22568_n8944 0.934191f
C3970 a_40396_n3237 VDD 0.338239f
C3971 a_31961_1204 VDD 0.490365f
C3972 a_45236_n9412 a_45684_n9412 0.013276f
C3973 a_25685_n7463 VDD 0.538324f
C3974 a_22772_n10512 VDD 0.299818f
C3975 a_36724_n12548 a_37172_n12548 0.013276f
C3976 a_45772_n12645 a_46132_n12548 0.087066f
C3977 a_47028_n12548 VDD 0.206217f
C3978 a_41740_n14213 a_42100_n14116 0.087066f
C3979 a_32308_n1976 a_35288_n1975 0.484997f
C3980 a_47028_n15684 VDD 0.206217f
C3981 a_45772_n15781 a_45684_n15684 0.285629f
C3982 a_36948_n15684 a_37396_n15684 0.013276f
C3983 a_44004_n1192 a_45100_1467 0.031635f
C3984 a_28212_n18820 VDD 0.205948f
C3985 a_28144_n4708 a_30740_n7464 0.381094f
C3986 a_41740_n4805 a_42100_n4708 0.087066f
C3987 a_47564_n4805 a_48012_n4805 0.012882f
C3988 a_46668_n17349 a_47028_n17252 0.087066f
C3989 a_47564_n101 VDD 0.312443f
C3990 a_44876_n18917 a_45324_n18917 0.012882f
C3991 a_31436_n18917 a_31796_n18820 0.087066f
C3992 a_24264_n6976 a_24576_n6976 0.119687f
C3993 a_24233_n3980 VDD 0.506821f
C3994 a_27281_n16854 a_27391_n11384 0.061428f
C3995 a_24041_816 VDD 0.261872f
C3996 a_44452_n7464 VDD 0.220197f
C3997 a_42300_n15348 CLK 0.048577f
C3998 a_42212_n10600 VDD 0.206217f
C3999 a_22600_n12124 a_22052_n15304 0.015199f
C4000 a_35604_n13736 VDD 0.208855f
C4001 a_43892_n14116 a_44340_n14116 0.013276f
C4002 a_31324_n4372 a_31656_n704 0.068873f
C4003 a_34012_n16916 VDD 0.315469f
C4004 a_48012_n3237 a_47924_n3140 0.285629f
C4005 a_43444_n3140 a_43892_n3140 0.013276f
C4006 a_33588_n3461 a_33416_n4240 0.011422f
C4007 a_24631_n3588 a_29560_n3544 0.028185f
C4008 a_21604_n20008 VDD 0.221763f
C4009 a_41204_1243 a_43833_1204 0.019043f
C4010 a_41616_1564 a_41864_1394 0.354223f
C4011 a_30676_n17252 a_30788_n18440 0.026657f
C4012 a_47028_n17252 a_47476_n17252 0.013276f
C4013 a_23479_n5156 a_22968_n6679 0.010442f
C4014 a_22444_n5156 a_21812_n6643 0.05004f
C4015 a_24492_n5156 a_28644_n9815 0.032173f
C4016 a_42636_n18917 a_42548_n18820 0.285629f
C4017 a_30408_n1104 VDD 0.369696f
C4018 a_38268_n20485 a_38716_n20485 0.013103f
C4019 a_26396_n20485 a_26308_n20388 0.285629f
C4020 a_29532_n10311 a_29992_n11150 0.0558f
C4021 a_32732_n10556 a_32628_n10512 0.026665f
C4022 a_28972_n7819 VDD 0.011991f
C4023 a_30787_n12167 a_30599_n12167 0.247613f
C4024 a_40308_n12548 a_40420_n13736 0.026657f
C4025 a_46020_n13736 VDD 0.210736f
C4026 a_46916_n1572 a_47364_n1572 0.013276f
C4027 a_38740_n14116 a_38628_n15304 0.026657f
C4028 a_44004_n1192 a_43556_n661 0.195747f
C4029 a_47812_n16872 VDD 0.211703f
C4030 a_22568_n4240 a_22772_n4240 0.66083f
C4031 a_30788_n16872 a_31236_n16872 0.013276f
C4032 a_23136_447 a_24913_864 0.153996f
C4033 a_35268_n20008 VDD 0.206217f
C4034 a_28436_n18440 a_28076_n18484 0.086905f
C4035 a_37844_n17252 a_37732_n18440 0.026657f
C4036 a_41764_n7464 a_41404_n7508 0.087066f
C4037 a_39636_n18820 a_40084_n18820 0.013276f
C4038 a_30396_n7508 a_28764_n8247 0.012963f
C4039 a_46556_n1236 VDD 0.299954f
C4040 a_25573_n12167 a_22220_n12996 0.995721f
C4041 a_41852_n9076 a_42300_n9076 0.012882f
C4042 a_38716_n20485 a_38628_n20388 0.285629f
C4043 a_23228_n6679 VDD 0.299057f
C4044 a_39524_n10600 a_39164_n10644 0.087066f
C4045 a_28456_n364 a_30781_n452 0.014892f
C4046 a_40308_n7844 VDD 0.212323f
C4047 a_26563_n12212 a_26239_n12996 0.016345f
C4048 a_41764_n12168 a_42212_n12168 0.013276f
C4049 a_37732_n12168 a_37820_n12212 0.285629f
C4050 a_47564_n11077 VDD 0.315469f
C4051 a_34708_n13736 a_34796_n13780 0.285629f
C4052 a_47476_n12548 a_47364_n13736 0.026657f
C4053 a_22600_n12124 a_22588_n15781 0.030975f
C4054 a_30372_376 a_30781_n452 0.018066f
C4055 a_38380_n14213 VDD 0.343298f
C4056 a_36500_n15304 a_36140_n15348 0.086635f
C4057 a_33004_n15348 a_33452_n15348 0.013103f
C4058 a_45684_n14116 a_45572_n15304 0.026657f
C4059 a_26499_n2732 a_27348_n2672 0.068207f
C4060 a_45324_n17349 VDD 0.324845f
C4061 a_46132_n3140 a_46020_n4328 0.026657f
C4062 a_32359_n4372 a_33015_n4284 0.510371f
C4063 a_41404_n20052 VDD 0.328902f
C4064 a_22444_n5156 a_32560_n7020 0.118346f
C4065 a_35716_n18440 a_36164_n18440 0.013276f
C4066 a_22264_n5852 a_23619_n6724 0.214675f
C4067 a_32132_n18440 a_32220_n18484 0.285629f
C4068 a_45212_n7508 a_45660_n7508 0.012552f
C4069 a_32692_n18820 a_32580_n20008 0.026657f
C4070 a_46916_n7464 a_47004_n7508 0.285629f
C4071 a_32308_n1976 VDD 0.290295f
C4072 a_23619_n9860 a_22264_n10556 0.226364f
C4073 a_38628_n20388 a_39076_n20388 0.013276f
C4074 a_35940_2475 OUT[2] 0.010684f
C4075 a_46668_n4805 VDD 0.318039f
C4076 a_46020_n10600 a_46468_n10600 0.013276f
C4077 a_25020_n11383 a_26563_n12212 0.06466f
C4078 a_28617_n8548 VDD 0.325011f
C4079 a_31760_n12168 a_31789_n12996 0.046256f
C4080 a_26431_n12168 VDD 0.699099f
C4081 a_43556_n13736 a_44004_n13736 0.013276f
C4082 a_39972_n13736 a_40060_n13780 0.285629f
C4083 a_42996_n14116 VDD 0.205948f
C4084 a_34649_n2412 a_34544_n2272 0.119281f
C4085 a_40420_n15304 a_40060_n15348 0.087066f
C4086 a_22500_n1976 a_22820_n2804 0.010732f
C4087 a_30104_n1148 a_29856_n1121 0.343084f
C4088 a_46132_n17252 VDD 0.210512f
C4089 a_41764_n16872 a_41852_n16916 0.285629f
C4090 a_37820_n16916 a_38268_n16916 0.012882f
C4091 a_41764_n4328 a_41852_n4372 0.285629f
C4092 a_37372_n20485 VDD 0.302862f
C4093 a_45124_n5896 a_45212_n5940 0.285629f
C4094 a_46468_n5896 a_46916_n5896 0.013276f
C4095 a_25276_n20052 a_25724_n20052 0.012882f
C4096 a_39636_n18820 a_39524_n20008 0.026657f
C4097 a_46020_n1572 VDD 0.207964f
C4098 a_28624_n9394 a_30472_n9815 0.012865f
C4099 a_22772_n5808 VDD 0.299581f
C4100 a_41852_n13780 CLK 0.013107f
C4101 a_27281_n16854 a_25831_n12996 0.352769f
C4102 a_24964_n14116 a_28121_n10980 0.660833f
C4103 a_40956_n9076 VDD 0.330158f
C4104 a_28300_n15348 a_31960_n13648 0.02824f
C4105 a_40868_n12168 VDD 0.208618f
C4106 a_22600_n12124 a_22588_n16916 0.012923f
C4107 a_36140_n13780 a_36140_n14213 0.05841f
C4108 a_45572_n13736 a_45212_n13780 0.086905f
C4109 a_46916_n15304 a_47364_n15304 0.013276f
C4110 a_44228_n2760 a_44316_n2804 0.285629f
C4111 a_45572_n15304 a_45660_n15348 0.285629f
C4112 a_40652_n1572 a_41684_n1976 0.023977f
C4113 a_34820_n18440 VDD 0.206217f
C4114 a_45212_n4372 a_45660_n4372 0.012552f
C4115 a_47364_n16872 a_47004_n16916 0.086742f
C4116 a_46916_n4328 a_47004_n4372 0.285629f
C4117 a_40260_n408 a_39804_464 0.024417f
C4118 a_37732_n20388 VDD 0.21066f
C4119 a_25612_n6679 a_25972_n6276 0.107156f
C4120 a_41852_n18484 a_42300_n18484 0.012882f
C4121 a_44428_n7941 a_44876_n7941 0.012882f
C4122 a_37260_n7941 a_37620_n7844 0.087174f
C4123 a_46580_n18820 a_46468_n20008 0.026657f
C4124 a_32580_n20008 a_32220_n20052 0.087066f
C4125 a_34649_n2412 VDD 0.986409f
C4126 a_29532_n10311 a_30296_n10980 0.046097f
C4127 a_45572_n5896 VDD 0.213324f
C4128 a_37484_n11077 a_37932_n11077 0.013103f
C4129 a_30871_n11728 a_30787_n12167 0.511257f
C4130 a_27281_n16854 VDD 1.19617f
C4131 a_22264_n13692 VDD 0.39292f
C4132 a_33077_n1191 a_32636_n2020 0.018292f
C4133 a_43196_n13780 a_43084_n14213 0.026339f
C4134 a_46020_n15304 VDD 0.210736f
C4135 a_22164_n2760 a_22876_n4284 0.048664f
C4136 a_40956_n18484 VDD 0.330158f
C4137 a_23564_n20836 a_24380_n18917 0.012909f
C4138 a_23207_n4708 a_22564_n5112 0.021488f
C4139 a_42748_n4372 a_42636_n4805 0.026339f
C4140 a_35244_n17349 a_35692_n17349 0.012882f
C4141 a_25530_n5112 a_24180_n5112 0.015598f
C4142 a_42636_n6373 a_43084_n6373 0.012882f
C4143 a_30808_n6334 a_31936_n6592 0.048436f
C4144 a_39076_n20008 a_39524_n20008 0.013276f
C4145 a_47452_n2804 VDD 0.313885f
C4146 a_42188_n9509 a_42100_n9412 0.285629f
C4147 a_22220_n12996 a_26531_n10207 0.020576f
C4148 a_41740_n6373 VDD 0.328902f
C4149 a_40620_n11077 a_40532_n10980 0.285629f
C4150 a_42100_n17252 CLK 0.020589f
C4151 a_34572_n12645 a_34932_n12548 0.087174f
C4152 a_43532_n12645 a_43980_n12645 0.012882f
C4153 a_22264_n13692 a_21604_n13252 0.1001f
C4154 a_42636_n12645 VDD 0.313885f
C4155 a_21772_n12996 a_23396_n16872 0.011036f
C4156 a_42188_n15781 VDD 0.313885f
C4157 a_33588_n3461 a_34348_n3140 0.011851f
C4158 a_34796_n15781 a_34708_n15684 0.285629f
C4159 a_43084_n15781 a_43532_n15781 0.012882f
C4160 a_32780_n18917 VDD 0.347953f
C4161 a_35692_n17349 a_36052_n17252 0.087066f
C4162 a_33900_n18917 a_34348_n18917 0.012882f
C4163 a_30740_n7464 a_30396_n7508 0.039324f
C4164 a_22264_n8988 a_22568_n8944 0.01851f
C4165 a_29532_n10311 a_33832_n8572 0.024738f
C4166 a_39948_n3237 VDD 0.330941f
C4167 a_31544_1248 VDD 1.34912f
C4168 a_24264_n6976 VDD 1.366f
C4169 a_43444_n10980 a_43892_n10980 0.013276f
C4170 a_24128_n10112 VDD 0.026027f
C4171 a_45772_n12645 a_45684_n12548 0.285629f
C4172 a_46580_n12548 VDD 0.209016f
C4173 a_32308_n1976 a_34223_n1976 0.021452f
C4174 a_41740_n14213 a_41652_n14116 0.285629f
C4175 a_46580_n15684 VDD 0.209016f
C4176 a_45324_n15781 a_45684_n15684 0.087066f
C4177 a_41292_n3237 a_41740_n3237 0.012882f
C4178 a_44004_n1192 a_43728_1248 0.029586f
C4179 a_27764_n18820 VDD 0.206173f
C4180 a_28144_n4708 a_31068_n6276 0.012484f
C4181 a_41740_n4805 a_41652_n4708 0.285629f
C4182 a_46668_n17349 a_46580_n17252 0.285629f
C4183 a_36052_n17252 a_36500_n17252 0.013276f
C4184 a_47116_n101 VDD 0.312206f
C4185 a_31436_n18917 a_31348_n18820 0.285629f
C4186 a_24681_n7116 a_24576_n6976 0.116059f
C4187 a_26095_n7464 a_26719_n7464 0.104193f
C4188 a_25948_n20485 a_26396_n20485 0.012552f
C4189 a_21872_n9394 a_25831_n11428 0.092815f
C4190 a_23404_816 VDD 0.485336f
C4191 a_27281_n16854 a_27167_n10808 0.031028f
C4192 a_38740_n9412 a_38628_n10600 0.026657f
C4193 a_41852_n15348 CLK 0.013107f
C4194 a_44004_n7464 VDD 0.21095f
C4195 a_23564_n11428 a_25132_n16432 0.488494f
C4196 a_37396_n10980 a_37284_n12168 0.026657f
C4197 a_23564_n8292 a_24752_n16132 0.304249f
C4198 a_41764_n10600 VDD 0.206217f
C4199 a_47476_n12548 a_47924_n12548 0.013276f
C4200 a_35156_n13736 VDD 0.208855f
C4201 a_27820_n16432 a_23564_n17700 0.036865f
C4202 a_46556_n1669 a_47004_n1669 0.012222f
C4203 a_33564_n16916 VDD 0.315469f
C4204 a_33812_n15684 a_33924_n16872 0.026657f
C4205 a_47476_n15684 a_47924_n15684 0.013276f
C4206 a_47564_n3237 a_47924_n3140 0.087066f
C4207 a_41204_1243 a_43416_1248 0.042802f
C4208 a_29332_1243 a_28492_332 0.037364f
C4209 a_46132_n4708 a_46580_n4708 0.013276f
C4210 a_22544_n4690 a_23619_n6724 0.02868f
C4211 a_28660_n18820 a_29108_n18820 0.013276f
C4212 a_42188_n18917 a_42548_n18820 0.087066f
C4213 a_45684_n6276 a_45572_n7464 0.026657f
C4214 a_23479_n5156 a_25724_n14564 0.033923f
C4215 a_30204_n1104 VDD 0.010384f
C4216 a_22264_n8988 a_22264_n10556 0.051236f
C4217 a_39076_n9032 a_39524_n9032 0.013276f
C4218 a_25948_n20485 a_26308_n20388 0.086905f
C4219 a_29532_n10311 a_25724_n14564 0.394457f
C4220 a_44452_n4328 VDD 0.220197f
C4221 a_45684_n9412 a_45572_n10600 0.026657f
C4222 a_34089_n10252 a_35392_n10172 0.01206f
C4223 a_28927_n10160 a_29479_n13735 0.104402f
C4224 a_45572_n13736 VDD 0.213324f
C4225 a_25577_n14956 a_25160_n14816 0.633318f
C4226 a_24220_n15260 a_24116_n15216 0.026665f
C4227 a_22500_n1976 a_22588_n2020 0.273845f
C4228 a_47364_n16872 VDD 0.205948f
C4229 a_41204_n15684 a_41316_n16872 0.026657f
C4230 a_34820_n20008 VDD 0.206217f
C4231 a_23728_464 a_23524_464 0.068207f
C4232 a_27988_n18440 a_28076_n18484 0.285629f
C4233 a_23932_n18484 a_24380_n18484 0.013103f
C4234 a_41316_n7464 a_41404_n7508 0.285629f
C4235 a_37372_n7508 a_37820_n7508 0.012882f
C4236 a_25524_n18820 a_25636_n20008 0.026657f
C4237 a_46108_n1236 VDD 0.300599f
C4238 a_25860_n20388 a_26308_n20388 0.013276f
C4239 a_38268_n20485 a_38628_n20388 0.087174f
C4240 a_23207_n4708 VDD 1.02114f
C4241 a_42548_n12548 CLK 0.029747f
C4242 a_39076_n10600 a_39164_n10644 0.285629f
C4243 a_26239_n11428 a_25559_n10980 0.15296f
C4244 a_42660_n10600 a_43108_n10600 0.013276f
C4245 a_28456_n364 a_28352_n320 0.084381f
C4246 a_39860_n7844 VDD 0.209112f
C4247 a_42548_n15684 CLK 0.029747f
C4248 a_37732_n12168 a_37372_n12212 0.087066f
C4249 a_23564_n11428 a_23816_n13248 0.015042f
C4250 a_26563_n12212 a_25831_n12996 0.026794f
C4251 a_47116_n11077 VDD 0.315469f
C4252 a_22600_n12124 a_22140_n15781 0.029702f
C4253 a_36052_n13736 a_36500_n13736 0.013276f
C4254 a_22876_n1148 a_23816_n704 0.056721f
C4255 a_24631_n3588 a_30451_n452 0.024354f
C4256 a_37932_n14213 VDD 0.328074f
C4257 a_36052_n15304 a_36140_n15348 0.285629f
C4258 a_27452_n2716 a_28454_n2424 0.035978f
C4259 a_27988_n4328 a_27337_n3140 0.075257f
C4260 a_44876_n17349 VDD 0.360805f
C4261 a_34460_n16916 a_34908_n16916 0.012552f
C4262 a_32359_n4372 a_33120_n3884 0.042802f
C4263 a_31787_n3969 a_33015_n4284 0.020455f
C4264 a_40956_n20052 VDD 0.328902f
C4265 a_28492_332 a_31076_376 0.721549f
C4266 a_32132_n18440 a_31772_n18484 0.087066f
C4267 a_41876_n5896 a_42324_n5896 0.013276f
C4268 a_22264_n5852 a_22968_n6679 0.187988f
C4269 a_22052_n20008 a_22500_n20008 0.013276f
C4270 a_46916_n7464 a_46556_n7508 0.086742f
C4271 a_24492_n5156 a_29444_n10116 0.04663f
C4272 a_29532_n10311 a_31460_n10116 0.010568f
C4273 a_46220_n4805 VDD 0.31977f
C4274 a_43644_n12212 a_44092_n12212 0.012882f
C4275 a_26563_n12212 VDD 0.442928f
C4276 a_39972_n13736 a_39612_n13780 0.087066f
C4277 a_42548_n14116 VDD 0.205948f
C4278 a_39972_n15304 a_40060_n15348 0.285629f
C4279 a_43556_n15304 a_44004_n15304 0.013276f
C4280 a_45684_n17252 VDD 0.212747f
C4281 a_41764_n4328 a_41404_n4372 0.087174f
C4282 a_41764_n16872 a_41404_n16916 0.087066f
C4283 a_36924_n20485 VDD 0.338856f
C4284 a_23484_n18484 a_23484_n18917 0.05841f
C4285 a_38628_n18440 a_39076_n18440 0.013276f
C4286 a_45572_n1572 VDD 0.208696f
C4287 a_24128_n5408 VDD 0.025152f
C4288 a_41852_n10644 a_41740_n11077 0.026339f
C4289 a_25559_n10980 a_24684_n16432 0.239204f
C4290 a_40508_n9076 VDD 0.313885f
C4291 a_38268_n12212 a_38156_n12645 0.026339f
C4292 a_40420_n12168 VDD 0.205948f
C4293 a_45124_n13736 a_45212_n13780 0.285629f
C4294 a_46468_n13736 a_46916_n13736 0.013276f
C4295 a_27988_n20388 VDD 1.79245f
C4296 a_22820_n2804 a_22052_n4708 0.015829f
C4297 a_27628_n3841 a_27337_n3140 0.309651f
C4298 a_45572_n15304 a_45212_n15348 0.086905f
C4299 a_44228_n2760 a_43868_n2804 0.086635f
C4300 a_40652_n1572 a_41292_n1669 0.017975f
C4301 a_34372_n18440 VDD 0.206217f
C4302 a_46916_n4328 a_46556_n4372 0.086742f
C4303 a_45212_n16916 a_45660_n16916 0.012552f
C4304 a_46916_n16872 a_47004_n16916 0.285629f
C4305 a_47028_n4 VDD 0.207033f
C4306 a_37284_n20388 VDD 0.208438f
C4307 a_30876_n18484 a_30988_n18917 0.026339f
C4308 a_32132_n20008 a_32220_n20052 0.285629f
C4309 a_35716_n20008 a_36164_n20008 0.013276f
C4310 a_37260_n7941 a_37172_n7844 0.285629f
C4311 a_38380_n9509 a_38828_n9509 0.013103f
C4312 a_45124_n5896 VDD 0.264203f
C4313 a_47452_n12212 a_47564_n12645 0.026339f
C4314 a_47004_n1236 a_47452_n1236 0.012222f
C4315 a_45572_n15304 VDD 0.213324f
C4316 a_31324_n4372 a_25084_1564 0.042005f
C4317 a_40508_n18484 VDD 0.313885f
C4318 a_25237_n5895 a_24180_n5112 0.010465f
C4319 a_23564_n20836 a_23932_n18917 0.048088f
C4320 a_45660_n16916 a_45772_n17349 0.026339f
C4321 a_30215_n6265 a_31936_n6592 0.401636f
C4322 a_37820_n18484 a_37932_n18917 0.026339f
C4323 a_22588_n18917 a_23036_n18917 0.013103f
C4324 a_41204_n7844 a_41652_n7844 0.013276f
C4325 a_47004_n2804 VDD 0.313885f
C4326 a_41740_n9509 a_42100_n9412 0.087066f
C4327 a_28736_1944 VDD 0.56452f
C4328 a_41292_n6373 VDD 0.335119f
C4329 a_24964_n14116 a_28009_n12168 0.029182f
C4330 a_40172_n11077 a_40532_n10980 0.086742f
C4331 a_48012_n9509 VDD 0.343411f
C4332 a_34572_n12645 a_34484_n12548 0.285629f
C4333 a_42188_n12645 VDD 0.313885f
C4334 a_35849_n1192 a_35916_n4 0.02049f
C4335 a_38828_n14213 a_39276_n14213 0.012882f
C4336 a_21772_n12996 a_22948_n16872 0.011877f
C4337 a_42972_n1236 a_42244_n1572 0.031722f
C4338 a_41740_n15781 VDD 0.313885f
C4339 a_33588_n3461 a_34860_n3189 0.05539f
C4340 a_25237_n4327 a_22052_n4708 0.06231f
C4341 a_34348_n15781 a_34708_n15684 0.087066f
C4342 a_24631_n3588 a_27452_n2716 0.048133f
C4343 a_25084_1564 a_31961_1204 0.02252f
C4344 a_32332_n18917 VDD 0.321441f
C4345 a_45772_n17349 a_46220_n17349 0.012882f
C4346 a_35692_n17349 a_35604_n17252 0.285629f
C4347 a_48012_n6373 a_47924_n6276 0.285629f
C4348 a_24492_n5156 a_28225_n9031 0.100639f
C4349 a_47004_n18484 a_47116_n18917 0.026339f
C4350 a_42548_n6276 a_42996_n6276 0.013276f
C4351 a_41852_n20052 a_42300_n20052 0.012882f
C4352 a_33116_n20052 a_33116_n20485 0.05841f
C4353 a_22016_n8961 a_22568_n8944 0.361958f
C4354 a_22264_n8988 a_22364_n8944 0.106759f
C4355 a_39500_n3237 VDD 0.320901f
C4356 a_32581_n9860 a_32628_n10512 0.01349f
C4357 a_44788_n9412 a_45236_n9412 0.013276f
C4358 a_30500_1564 VDD 0.302073f
C4359 a_24681_n7116 VDD 0.495192f
C4360 a_45324_n12645 a_45684_n12548 0.087066f
C4361 a_36276_n12548 a_36724_n12548 0.013276f
C4362 a_46132_n12548 VDD 0.210512f
C4363 a_41292_n14213 a_41652_n14116 0.087066f
C4364 a_32308_n1976 a_33999_n1400 0.022666f
C4365 a_46132_n15684 VDD 0.210512f
C4366 a_36500_n15684 a_36948_n15684 0.013276f
C4367 a_45324_n15781 a_45236_n15684 0.285629f
C4368 a_27316_n18820 VDD 0.206648f
C4369 a_44004_n1192 a_43833_1204 0.065966f
C4370 a_46220_n17349 a_46580_n17252 0.087066f
C4371 a_27988_n4328 a_25831_n11428 0.036748f
C4372 a_41292_n4805 a_41652_n4708 0.087066f
C4373 a_47116_n4805 a_47564_n4805 0.012882f
C4374 a_46668_n101 VDD 0.314754f
C4375 a_30988_n18917 a_31348_n18820 0.087066f
C4376 a_44428_n18917 a_44876_n18917 0.012882f
C4377 a_25685_n7463 a_26719_n7464 0.054912f
C4378 a_40060_n20052 a_40060_n20485 0.05841f
C4379 a_27485_n8500 a_25831_n11428 0.014596f
C4380 a_23136_447 VDD 1.0648f
C4381 a_43556_n7464 VDD 0.209375f
C4382 a_27055_n12168 a_27279_n12146 0.538085f
C4383 a_23564_n8292 a_24088_n16087 0.246759f
C4384 a_24569_n11820 a_25880_n11708 0.010064f
C4385 a_26547_n12951 a_26983_n12728 0.015613f
C4386 a_24964_n14116 a_27744_n12908 0.04904f
C4387 a_41316_n10600 VDD 0.206217f
C4388 a_34708_n13736 VDD 0.13106f
C4389 a_43444_n14116 a_43892_n14116 0.013276f
C4390 a_33116_n16916 VDD 0.332191f
C4391 a_42996_n3140 a_43444_n3140 0.013276f
C4392 a_47564_n3237 a_47476_n3140 0.285629f
C4393 a_22544_n4690 a_22968_n6679 0.048728f
C4394 a_46580_n17252 a_47028_n17252 0.013276f
C4395 a_30228_n17252 a_30340_n18440 0.026657f
C4396 a_33048_n7420 a_34176_n6976 0.048436f
C4397 a_24672_n11339 a_22220_n12996 0.036211f
C4398 a_32856_n7376 a_33497_n9032 0.022479f
C4399 a_42188_n18917 a_42100_n18820 0.285629f
C4400 a_30716_n1148 VDD 0.267951f
C4401 a_25948_n20485 a_25860_n20388 0.285629f
C4402 a_37820_n20485 a_38268_n20485 0.013103f
C4403 a_44004_n4328 VDD 0.2115f
C4404 a_34089_n10252 a_33672_n10112 0.633318f
C4405 a_30576_376 VDD 0.010406f
C4406 a_30787_n12167 a_31760_n12168 0.484748f
C4407 a_39860_n12548 a_39972_n13736 0.026657f
C4408 a_45124_n13736 VDD 0.26277f
C4409 a_38292_n14116 a_38180_n15304 0.026657f
C4410 a_46468_n1572 a_46916_n1572 0.013276f
C4411 a_46916_n16872 VDD 0.205962f
C4412 a_30340_n16872 a_30788_n16872 0.013276f
C4413 a_22876_n4284 a_22772_n4240 0.026665f
C4414 a_22116_860 a_22340_376 0.013419f
C4415 a_34372_n20008 VDD 0.206217f
C4416 a_37396_n17252 a_37284_n18440 0.026657f
C4417 a_27988_n18440 a_27628_n18484 0.086905f
C4418 a_39188_n18820 a_39636_n18820 0.013276f
C4419 a_41316_n7464 a_40956_n7508 0.087066f
C4420 a_45660_n1236 VDD 0.303781f
C4421 a_25831_n11428 a_26470_n9322 0.03648f
C4422 a_41404_n9076 a_41852_n9076 0.012882f
C4423 a_28617_n8548 a_30472_n9815 0.483776f
C4424 a_38268_n20485 a_38180_n20388 0.285629f
C4425 a_26358_n4618 VDD 0.759349f
C4426 a_42100_n12548 CLK 0.020589f
C4427 a_48012_332 VDD 0.324628f
C4428 a_39076_n10600 a_38716_n10644 0.087066f
C4429 a_28456_n364 a_30451_n452 0.212448f
C4430 a_39412_n7844 VDD 0.210723f
C4431 a_42100_n15684 CLK 0.020589f
C4432 a_23564_n11428 a_24233_n13388 0.011641f
C4433 a_37284_n12168 a_37372_n12212 0.285629f
C4434 a_41316_n12168 a_41764_n12168 0.013276f
C4435 a_46668_n11077 VDD 0.318039f
C4436 a_47028_n12548 a_46916_n13736 0.026657f
C4437 a_37484_n14213 VDD 0.322568f
C4438 a_45236_n14116 a_45124_n15304 0.026657f
C4439 a_36052_n15304 a_35692_n15348 0.087174f
C4440 a_28752_n15348 a_23564_n17700 0.016496f
C4441 a_44428_n17349 VDD 0.321554f
C4442 a_47924_n15684 a_47812_n16872 0.026657f
C4443 a_31787_n3969 a_33120_n3884 0.019033f
C4444 a_45684_n3140 a_45572_n4328 0.026657f
C4445 a_30372_376 a_24631_n3588 0.038899f
C4446 a_40508_n20052 VDD 0.328237f
C4447 a_22444_n5156 a_31799_n7508 0.010538f
C4448 a_31684_n18440 a_31772_n18484 0.285629f
C4449 a_21604_n5412 a_23619_n6724 0.030097f
C4450 a_35268_n18440 a_35716_n18440 0.013276f
C4451 a_32244_n18820 a_32132_n20008 0.026657f
C4452 a_46468_n7464 a_46556_n7508 0.285629f
C4453 a_38180_n20388 a_38628_n20388 0.013276f
C4454 a_29532_n10311 a_30136_n10600 0.042947f
C4455 a_45772_n4805 VDD 0.321879f
C4456 a_30871_n11728 a_34350_n10980 0.072763f
C4457 a_45572_n10600 a_46020_n10600 0.013276f
C4458 a_24152_n11680 VDD 1.36876f
C4459 a_39524_n13736 a_39612_n13780 0.285629f
C4460 a_43108_n13736 a_43556_n13736 0.013276f
C4461 a_30716_n1148 a_31656_n704 0.056721f
C4462 VDD OUT[2] 0.965382f
C4463 a_42100_n14116 VDD 0.205948f
C4464 a_39972_n15304 a_39612_n15348 0.087066f
C4465 a_30104_n1148 a_29444_n708 0.105951f
C4466 a_45236_n17252 VDD 0.229781f
C4467 a_41316_n16872 a_41404_n16916 0.285629f
C4468 a_37372_n16916 a_37820_n16916 0.012882f
C4469 a_26271_n4306 a_26358_n4618 0.018499f
C4470 a_41316_n4328 a_41404_n4372 0.285629f
C4471 a_36252_n20485 VDD 0.325169f
C4472 a_23404_816 a_24628_n363 0.017885f
C4473 a_46020_n5896 a_46468_n5896 0.013276f
C4474 a_28772_n20008 a_28860_n20052 0.285629f
C4475 a_39188_n18820 a_39076_n20008 0.026657f
C4476 a_24828_n20052 a_25276_n20052 0.012882f
C4477 a_45124_n1572 VDD 0.232927f
C4478 a_29800_n9815 a_28624_n9394 0.516665f
C4479 a_40060_n9076 VDD 0.314419f
C4480 a_42748_n16916 CLK 0.012909f
C4481 a_23949_n12996 a_24573_n12996 0.104193f
C4482 a_28300_n15348 a_31455_n13648 0.01218f
C4483 a_39972_n12168 VDD 0.207295f
C4484 a_35692_n13780 a_35692_n14213 0.05841f
C4485 a_45124_n15304 a_45212_n15348 0.285629f
C4486 a_43780_n2760 a_43868_n2804 0.285629f
C4487 a_46468_n15304 a_46916_n15304 0.013276f
C4488 a_40652_n1572 a_40196_n1884 0.286545f
C4489 a_33924_n18440 VDD 0.206217f
C4490 a_46916_n16872 a_46556_n16916 0.086742f
C4491 a_46468_n4328 a_46556_n4372 0.285629f
C4492 a_22052_n4708 a_36773_n5468 0.01135f
C4493 a_36836_n20388 VDD 0.227486f
C4494 a_41404_n18484 a_41852_n18484 0.012882f
C4495 a_24492_n5156 a_28121_n10980 0.020187f
C4496 a_46132_n18820 a_46020_n20008 0.026657f
C4497 a_43980_n7941 a_44428_n7941 0.012882f
C4498 a_36812_n7941 a_37172_n7844 0.087174f
C4499 a_32132_n20008 a_31772_n20052 0.087066f
C4500 a_42636_n11077 CLK 0.01698f
C4501 a_27281_n16854 a_28335_n10644 0.041627f
C4502 a_44204_n5940 VDD 0.356422f
C4503 a_24964_n14116 a_28300_n15348 0.15675f
C4504 a_37036_n11077 a_37484_n11077 0.013103f
C4505 a_21872_n12530 VDD 0.374448f
C4506 a_27496_n14116 a_27700_n14116 0.66083f
C4507 a_42748_n13780 a_42636_n14213 0.026339f
C4508 a_23004_n2332 a_26631_7 0.023677f
C4509 a_45124_n15304 VDD 0.26277f
C4510 a_22164_n2760 a_22016_n4257 0.044921f
C4511 a_40060_n18484 VDD 0.314419f
C4512 a_24672_n11339 a_24180_n5112 0.347613f
C4513 a_34796_n17349 a_35244_n17349 0.012882f
C4514 a_42300_n4372 a_42188_n4805 0.026339f
C4515 a_23564_n20836 a_23484_n18917 0.013207f
C4516 a_42188_n6373 a_42636_n6373 0.012882f
C4517 a_48012_n7941 a_47924_n7844 0.285629f
C4518 a_38628_n20008 a_39076_n20008 0.013276f
C4519 a_46556_n2804 VDD 0.31705f
C4520 a_22220_n12996 a_23816_n10112 0.010849f
C4521 a_22500_n1976 VDD 1.04209f
C4522 a_41740_n9509 a_41652_n9412 0.285629f
C4523 a_40396_n6373 VDD 0.349262f
C4524 a_40172_n11077 a_40084_n10980 0.285629f
C4525 a_23564_n8292 a_22948_n14820 0.013225f
C4526 a_47564_n9509 VDD 0.315469f
C4527 a_43084_n12645 a_43532_n12645 0.012882f
C4528 a_34124_n12645 a_34484_n12548 0.087174f
C4529 a_41740_n12645 VDD 0.313885f
C4530 a_21772_n12996 a_22500_n16872 0.014825f
C4531 a_41292_n15781 VDD 0.318502f
C4532 a_34348_n15781 a_34260_n15684 0.285629f
C4533 a_42636_n15781 a_43084_n15781 0.012882f
C4534 a_33588_n3461 a_34000_n3140 0.536965f
C4535 a_31884_n18917 VDD 0.323762f
C4536 a_31324_n4372 a_31856_1248 0.024258f
C4537 a_25084_1564 a_31544_1248 0.035966f
C4538 a_35244_n17349 a_35604_n17252 0.087066f
C4539 a_30320_n6636 a_31799_n7508 0.035221f
C4540 a_47564_n6373 a_47924_n6276 0.087066f
C4541 a_25612_n6679 a_33497_n9032 0.474841f
C4542 a_33452_n18917 a_33900_n18917 0.012882f
C4543 a_24492_n5156 a_29540_n11728 0.226646f
C4544 a_21604_n8548 a_22568_n8944 0.08126f
C4545 a_22016_n8961 a_22364_n8944 0.401636f
C4546 a_37585_n3140 VDD 0.554202f
C4547 a_30296_1564 VDD 0.368809f
C4548 a_42996_n10980 a_43444_n10980 0.013276f
C4549 a_27485_n10068 VDD 0.692579f
C4550 a_45324_n12645 a_45236_n12548 0.285629f
C4551 a_45684_n12548 VDD 0.212747f
C4552 a_41292_n14213 a_41204_n14116 0.285629f
C4553 a_45684_n15684 VDD 0.212747f
C4554 a_44876_n15781 a_45236_n15684 0.087066f
C4555 a_26868_n18820 VDD 0.206098f
C4556 a_31961_1204 a_31856_1248 0.116059f
C4557 a_44004_n1192 a_43416_1248 0.050588f
C4558 a_46220_n17349 a_46132_n17252 0.285629f
C4559 a_35604_n17252 a_36052_n17252 0.013276f
C4560 a_41292_n4805 a_41204_n4708 0.285629f
C4561 a_46220_n101 VDD 0.315647f
C4562 a_30988_n18917 a_30900_n18820 0.285629f
C4563 a_25685_n7463 a_26095_n7464 0.562529f
C4564 a_23016_n7376 a_23220_n7376 0.66083f
C4565 a_25500_n20485 a_25948_n20485 0.012552f
C4566 a_22568_n4240 VDD 0.362252f
C4567 a_38292_n9412 a_38180_n10600 0.026657f
C4568 a_22116_860 VDD 0.80662f
C4569 a_43108_n7464 VDD 0.206367f
C4570 a_24152_n11680 a_24464_n11680 0.119687f
C4571 a_26547_n12951 a_26635_n12996 0.124276f
C4572 a_24965_n9860 a_25844_n14116 0.017318f
C4573 a_40868_n10600 VDD 0.208618f
C4574 a_47028_n12548 a_47476_n12548 0.013276f
C4575 a_29479_n13735 VDD 0.963913f
C4576 a_46108_n1669 a_46556_n1669 0.013103f
C4577 a_31324_n4372 OUT[0] 0.028613f
C4578 a_32668_n16916 VDD 0.319553f
C4579 a_33364_n15684 a_33476_n16872 0.026657f
C4580 a_47116_n3237 a_47476_n3140 0.087066f
C4581 a_47028_n15684 a_47476_n15684 0.013276f
C4582 a_41204_1243 a_42168_1564 0.08126f
C4583 a_27736_1248 a_28132_376 0.022269f
C4584 a_45684_n4708 a_46132_n4708 0.013276f
C4585 a_28212_n18820 a_28660_n18820 0.013276f
C4586 a_32455_n7420 a_34176_n6976 0.401636f
C4587 a_45236_n6276 a_45124_n7464 0.026657f
C4588 a_41740_n18917 a_42100_n18820 0.087066f
C4589 a_29856_n1121 VDD 0.826427f
C4590 a_25500_n20485 a_25860_n20388 0.086905f
C4591 a_47564_n101 a_48012_n101 0.012001f
C4592 a_38628_n9032 a_39076_n9032 0.013276f
C4593 a_43556_n4328 VDD 0.209925f
C4594 a_25020_n11383 a_26543_n11384 0.035517f
C4595 a_45236_n9412 a_45124_n10600 0.026657f
C4596 a_44540_n13780 VDD 0.353322f
C4597 a_22500_n1976 a_21916_n1975 0.519844f
C4598 a_46468_n16872 VDD 0.209055f
C4599 a_24233_n3980 a_23816_n3840 0.633318f
C4600 a_24041_816 a_23728_464 0.386669f
C4601 a_33924_n20008 VDD 0.206217f
C4602 a_23404_816 a_23524_464 0.119099f
C4603 a_27540_n18440 a_27628_n18484 0.285629f
C4604 a_23484_n18484 a_23932_n18484 0.013103f
C4605 a_21812_n6643 a_24233_n8684 0.01496f
C4606 a_40868_n7464 a_40956_n7508 0.285629f
C4607 a_45212_n1236 VDD 0.325897f
C4608 a_37820_n20485 a_38180_n20388 0.087174f
C4609 a_25831_n11428 a_26266_n9240 0.029748f
C4610 a_28617_n8548 a_28624_n9394 0.076858f
C4611 a_25412_n20388 a_25860_n20388 0.013276f
C4612 a_25860_n9032 a_22220_n12996 0.02665f
C4613 a_26154_n4536 VDD 0.594685f
C4614 a_38628_n10600 a_38716_n10644 0.285629f
C4615 a_27281_n16854 a_27279_n12146 0.032786f
C4616 a_42212_n10600 a_42660_n10600 0.013276f
C4617 a_27485_n10068 a_27167_n10808 0.03239f
C4618 a_38964_n7844 VDD 0.212805f
C4619 a_46220_n11077 VDD 0.31977f
C4620 a_35604_n13736 a_36052_n13736 0.013276f
C4621 a_29812_860 a_30451_n452 0.028159f
C4622 a_37036_n14213 VDD 0.33541f
C4623 a_41204_n1572 a_41092_n2760 0.026657f
C4624 a_35604_n15304 a_35692_n15348 0.285629f
C4625 a_43980_n17349 VDD 0.31896f
C4626 a_34012_n16916 a_34460_n16916 0.012552f
C4627 a_40652_n1572 a_39308_n452 0.02788f
C4628 a_22052_n4708 a_22564_n5112 0.024906f
C4629 a_41864_1394 a_40260_n408 0.037788f
C4630 a_40060_n20052 VDD 0.297323f
C4631 a_41428_n5896 a_41876_n5896 0.013276f
C4632 a_21604_n5412 a_22968_n6679 0.032681f
C4633 a_31684_n18440 a_31324_n18484 0.087066f
C4634 a_22220_n9860 a_24264_n6976 0.033064f
C4635 a_21604_n20008 a_22052_n20008 0.013276f
C4636 a_24492_n5156 a_28435_n10599 0.024f
C4637 a_46468_n7464 a_46108_n7508 0.086905f
C4638 a_29532_n10311 a_29444_n10116 0.555195f
C4639 a_25573_n12167 a_25020_n11383 0.155f
C4640 a_45324_n4805 VDD 0.324845f
C4641 a_43196_n12212 a_43644_n12212 0.012882f
C4642 a_31760_n12168 a_31459_n12996 0.083495f
C4643 a_24569_n11820 VDD 0.504868f
C4644 a_39524_n13736 a_39164_n13780 0.087066f
C4645 a_35568_n4 a_35916_n4 0.401636f
C4646 a_29856_n1121 a_31656_n704 0.510371f
C4647 a_41652_n14116 VDD 0.205948f
C4648 a_43108_n15304 a_43556_n15304 0.013276f
C4649 a_39524_n15304 a_39612_n15348 0.285629f
C4650 a_44788_n17252 VDD 0.22479f
C4651 a_41316_n16872 a_40956_n16916 0.087066f
C4652 a_23564_n20836 a_24380_n18484 0.012909f
C4653 a_41316_n4328 a_40956_n4372 0.087174f
C4654 a_35804_n20485 VDD 0.296789f
C4655 a_23036_n18484 a_23036_n18917 0.05841f
C4656 a_38180_n18440 a_38628_n18440 0.013276f
C4657 a_28772_n20008 a_28412_n20052 0.086635f
C4658 a_31011_n8292 a_31341_n8292 0.538085f
C4659 a_44676_n1572 VDD 0.214954f
C4660 a_27281_n16854 a_28624_n9394 0.290765f
C4661 a_41404_n10644 a_41292_n11077 0.026339f
C4662 a_39612_n9076 VDD 0.317476f
C4663 a_42300_n16916 CLK 0.048577f
C4664 a_28300_n15348 a_32152_n13692 0.024725f
C4665 a_37820_n12212 a_37708_n12645 0.026339f
C4666 a_39524_n12168 VDD 0.209499f
C4667 a_46020_n13736 a_46468_n13736 0.013276f
C4668 a_43780_n2760 a_43420_n2804 0.087174f
C4669 a_40652_n1572 a_37221_n3543 0.04674f
C4670 a_33476_n18440 VDD 0.206217f
C4671 a_46468_n16872 a_46556_n16916 0.285629f
C4672 a_46468_n4328 a_46108_n4372 0.086905f
C4673 a_36164_n20388 VDD 0.209676f
C4674 a_30428_n18484 a_30540_n18917 0.026339f
C4675 a_25972_n6276 a_34392_n9815 0.526259f
C4676 a_36812_n7941 a_36724_n7844 0.285629f
C4677 a_35268_n20008 a_35716_n20008 0.013276f
C4678 a_31684_n20008 a_31772_n20052 0.285629f
C4679 a_32984_n2672 VDD 0.361102f
C4680 a_42188_n11077 CLK 0.047331f
C4681 a_37932_n9509 a_38380_n9509 0.013103f
C4682 a_43756_n5940 VDD 0.333483f
C4683 a_27526_n9816 VDD 0.326487f
C4684 a_31459_n12996 a_31789_n12996 0.538085f
C4685 a_47004_n12212 a_47116_n12645 0.026339f
C4686 a_23619_n12996 VDD 0.3147f
C4687 a_46556_n1236 a_47004_n1236 0.012222f
C4688 a_27804_n14165 a_28744_n14432 0.056721f
C4689 a_26944_n14116 a_29056_n14432 0.277491f
C4690 a_25844_n14116 a_25636_n14520 0.013419f
C4691 a_23004_n2332 a_26736_n364 0.017142f
C4692 a_44540_n15348 VDD 0.353322f
C4693 a_44540_n15348 a_44428_n15781 0.026339f
C4694 a_27085_n16132 a_27709_n16132 0.104193f
C4695 a_28736_1944 a_25084_1564 0.02084f
C4696 a_39612_n18484 VDD 0.317476f
C4697 a_45212_n16916 a_45324_n17349 0.026339f
C4698 a_37372_n18484 a_37484_n18917 0.026339f
C4699 a_22140_n18917 a_22588_n18917 0.013103f
C4700 a_47564_n7941 a_47924_n7844 0.087066f
C4701 a_22712_n7420 a_22220_n12996 0.022684f
C4702 a_46108_n2804 VDD 0.318654f
C4703 a_41292_n9509 a_41652_n9412 0.087066f
C4704 a_22220_n12996 a_24233_n10252 0.017217f
C4705 a_39948_n6373 VDD 0.329456f
C4706 a_39724_n11077 a_40084_n10980 0.086742f
C4707 a_47564_n11077 a_48012_n11077 0.012882f
C4708 a_47116_n9509 VDD 0.315469f
C4709 a_34124_n12645 a_34036_n12548 0.285629f
C4710 a_41292_n12645 VDD 0.320102f
C4711 a_21772_n12996 a_22052_n16872 0.054101f
C4712 a_38380_n14213 a_38828_n14213 0.012882f
C4713 a_40620_n15781 VDD 0.343849f
C4714 a_33900_n15781 a_34260_n15684 0.087066f
C4715 a_31324_n4372 a_31961_1204 0.011818f
C4716 a_25084_1564 a_30500_1564 0.014374f
C4717 a_31436_n18917 VDD 0.362787f
C4718 a_35244_n17349 a_35156_n17252 0.285629f
C4719 a_45324_n17349 a_45772_n17349 0.012882f
C4720 a_47564_n6373 a_47476_n6276 0.285629f
C4721 a_42100_n6276 a_42548_n6276 0.013276f
C4722 a_46556_n18484 a_46668_n18917 0.026339f
C4723 a_41404_n20052 a_41852_n20052 0.012882f
C4724 a_24492_n5156 a_28009_n12168 0.016679f
C4725 a_21604_n8548 a_22364_n8944 0.011851f
C4726 a_22016_n8961 a_22876_n8988 0.882105f
C4727 a_22052_n4708 VDD 1.37665f
C4728 a_44340_n9412 a_44788_n9412 0.013276f
C4729 a_30092_1564 VDD 0.01146f
C4730 a_26861_n10135 VDD 0.565226f
C4731 a_35828_n12548 a_36276_n12548 0.013276f
C4732 a_44876_n12645 a_45236_n12548 0.087066f
C4733 a_45236_n12548 VDD 0.229781f
C4734 a_32636_n2020 a_38312_n1975 0.194922f
C4735 a_40620_n14213 a_41204_n14116 0.016748f
C4736 a_45236_n15684 VDD 0.229781f
C4737 a_44876_n15781 a_44788_n15684 0.285629f
C4738 a_36052_n15684 a_36500_n15684 0.013276f
C4739 a_31544_1248 a_31856_1248 0.119687f
C4740 a_26420_n18820 VDD 0.206979f
C4741 a_46668_n4805 a_47116_n4805 0.012882f
C4742 a_40508_n4805 a_41204_n4708 0.012267f
C4743 a_45772_n17349 a_46132_n17252 0.087066f
C4744 a_28144_n4708 a_30808_n6334 0.015202f
C4745 a_24631_n3588 a_25612_n6679 0.043289f
C4746 a_45772_n101 VDD 0.321879f
C4747 a_43980_n18917 a_44428_n18917 0.012882f
C4748 a_30540_n18917 a_30900_n18820 0.087066f
C4749 a_39612_n20052 a_39612_n20485 0.05841f
C4750 a_22364_n4240 VDD 0.010384f
C4751 a_42660_n7464 VDD 0.206367f
C4752 a_26563_n12212 a_27279_n12146 0.053707f
C4753 a_26431_n12168 a_27055_n12168 0.104193f
C4754 a_24569_n11820 a_24464_n11680 0.116059f
C4755 a_26547_n12951 a_26239_n12996 0.118456f
C4756 a_24964_n14116 a_26635_n12996 0.019544f
C4757 a_40420_n10600 VDD 0.205948f
C4758 a_31960_n13648 VDD 0.251522f
C4759 a_42996_n14116 a_43444_n14116 0.013276f
C4760 a_32220_n16916 VDD 0.321588f
C4761 a_47116_n3237 a_47028_n3140 0.285629f
C4762 a_33588_n3461 a_33015_n4284 0.014454f
C4763 a_42548_n3140 a_42996_n3140 0.013276f
C4764 a_41204_1243 a_41964_1564 0.011851f
C4765 a_47924_n18820 VDD 0.213248f
C4766 a_29780_n17252 a_29892_n18440 0.026657f
C4767 a_46132_n17252 a_46580_n17252 0.013276f
C4768 a_32560_n7020 a_34176_n6976 0.011851f
C4769 a_41740_n18917 a_41652_n18820 0.285629f
C4770 a_24492_n5156 a_22220_n12996 0.037526f
C4771 a_22264_n8988 a_21772_n9860 0.026802f
C4772 a_25500_n20485 a_25412_n20388 0.285629f
C4773 a_37372_n20485 a_37820_n20485 0.013103f
C4774 a_45324_n101 a_45236_n4 0.285629f
C4775 a_43108_n4328 VDD 0.206917f
C4776 a_30808_n10116 a_30808_n10600 0.317701f
C4777 a_31872_n10529 a_33984_n10112 0.277491f
C4778 a_25020_n11383 a_26547_n12951 0.028183f
C4779 a_31011_n8292 VDD 0.340835f
C4780 a_26543_n11384 VDD 0.693087f
C4781 a_39412_n12548 a_39524_n13736 0.026657f
C4782 a_44092_n13780 VDD 0.3211f
C4783 a_23360_n15233 a_25472_n14816 0.277491f
C4784 a_46020_n1572 a_46468_n1572 0.013276f
C4785 a_37844_n14116 a_37732_n15304 0.026657f
C4786 a_46020_n16872 VDD 0.210736f
C4787 a_40532_n15684 a_40420_n16872 0.026657f
C4788 a_23136_447 a_23524_464 0.427756f
C4789 a_35849_n1192 a_35119_398 0.031814f
C4790 a_33476_n20008 VDD 0.206217f
C4791 a_27988_n4328 a_25724_n14564 0.030235f
C4792 a_27540_n18440 a_27180_n18484 0.086905f
C4793 a_38740_n18820 a_39188_n18820 0.013276f
C4794 a_40868_n7464 a_40508_n7508 0.087066f
C4795 a_24740_n18820 a_24740_n20008 0.05841f
C4796 a_47812_n1192 VDD 0.212403f
C4797 a_25831_n11428 a_25642_n9816 0.075958f
C4798 a_37820_n20485 a_37732_n20388 0.285629f
C4799 a_40956_n9076 a_41404_n9076 0.012882f
C4800 a_25530_n5112 VDD 0.799833f
C4801 a_27281_n16854 a_27055_n12168 0.013348f
C4802 a_25573_n12167 a_25831_n12996 0.123936f
C4803 a_38628_n10600 a_38268_n10644 0.087066f
C4804 a_38516_n7844 VDD 0.216736f
C4805 a_22600_n12124 a_21892_n12952 0.02569f
C4806 a_40868_n12168 a_41316_n12168 0.013276f
C4807 a_45772_n11077 VDD 0.321879f
C4808 a_22364_n1104 a_22568_n1104 0.048436f
C4809 a_22016_n1121 a_23816_n704 0.510371f
C4810 a_46580_n12548 a_46468_n13736 0.026657f
C4811 a_36588_n14213 VDD 0.299665f
C4812 a_35604_n15304 a_35244_n15348 0.087174f
C4813 a_31324_n4372 a_32308_n1976 0.016284f
C4814 a_43532_n17349 VDD 0.317216f
C4815 a_45236_n3140 a_45124_n4328 0.026657f
C4816 a_47476_n15684 a_47364_n16872 0.026657f
C4817 a_31787_n3969 a_32359_n4372 0.63615f
C4818 a_39612_n20052 VDD 0.30038f
C4819 a_29812_860 a_30372_376 0.302602f
C4820 a_34820_n18440 a_35268_n18440 0.013276f
C4821 a_31236_n18440 a_31324_n18484 0.285629f
C4822 a_22220_n9860 a_24681_n7116 0.022729f
C4823 a_37732_n5896 a_37820_n5940 0.285629f
C4824 a_46020_n7464 a_46108_n7508 0.285629f
C4825 a_31796_n18820 a_31684_n20008 0.026657f
C4826 a_47364_n7464 a_47812_n7464 0.013276f
C4827 a_37732_n20388 a_38180_n20388 0.013276f
C4828 a_44876_n4805 VDD 0.360805f
C4829 a_45124_n10600 a_45572_n10600 0.013276f
C4830 a_25573_n12167 VDD 1.45527f
C4831 a_35568_n4 a_36428_n53 0.882105f
C4832 a_29856_n1121 a_32073_n844 0.020455f
C4833 a_42660_n13736 a_43108_n13736 0.013276f
C4834 a_39076_n13736 a_39164_n13780 0.285629f
C4835 a_41204_n14116 VDD 0.226701f
C4836 a_37221_n3543 a_36217_n3500 0.111698f
C4837 a_34649_n2412 a_34232_n2272 0.612712f
C4838 a_39524_n15304 a_39164_n15348 0.087066f
C4839 a_44340_n17252 VDD 0.212126f
C4840 a_23564_n20836 a_23932_n18484 0.048002f
C4841 a_40868_n4328 a_40956_n4372 0.285629f
C4842 a_26047_n4328 a_26154_n4536 0.012528f
C4843 a_40868_n16872 a_40956_n16916 0.285629f
C4844 a_35356_n20485 VDD 0.296789f
C4845 a_29612_n8292 a_29123_n6679 0.337396f
C4846 a_45572_n5896 a_46020_n5896 0.013276f
C4847 a_38740_n18820 a_38628_n20008 0.026657f
C4848 a_24380_n20052 a_24828_n20052 0.012882f
C4849 a_28324_n20008 a_28412_n20052 0.285629f
C4850 a_44228_n1572 VDD 0.207706f
C4851 a_26470_n9322 a_25724_n14564 0.032965f
C4852 a_23816_n5408 VDD 1.35827f
C4853 a_26543_n11384 a_27167_n10808 0.104193f
C4854 a_41852_n16916 CLK 0.013107f
C4855 a_39164_n9076 VDD 0.319301f
C4856 a_28300_n15348 a_31559_n13692 0.064397f
C4857 a_22264_n13692 a_23949_n12996 0.018531f
C4858 a_21772_n12996 a_25831_n12996 0.390675f
C4859 a_39076_n12168 VDD 0.211414f
C4860 a_22600_n12124 a_23844_n16872 0.011176f
C4861 a_35244_n13780 a_35244_n14213 0.05841f
C4862 a_36500_n15304 VDD 0.21078f
C4863 a_46020_n15304 a_46468_n15304 0.013276f
C4864 a_43332_n2760 a_43420_n2804 0.285629f
C4865 a_33028_n18440 VDD 0.211234f
C4866 a_47364_n4328 a_47812_n4328 0.013276f
C4867 a_46020_n4328 a_46108_n4372 0.285629f
C4868 a_46468_n16872 a_46108_n16916 0.086905f
C4869 a_35716_n20388 VDD 0.203482f
C4870 a_40956_n18484 a_41404_n18484 0.012882f
C4871 a_31684_n20008 a_31324_n20052 0.087066f
C4872 a_45684_n18820 a_45572_n20008 0.026657f
C4873 a_43532_n7941 a_43980_n7941 0.012882f
C4874 a_36364_n7941 a_36724_n7844 0.087174f
C4875 a_32780_n2672 VDD 0.010618f
C4876 a_43308_n5940 VDD 0.331266f
C4877 a_36588_n11077 a_37036_n11077 0.013103f
C4878 a_27302_n9816 VDD 0.589121f
C4879 a_21772_n12996 VDD 1.46855f
C4880 a_26944_n14116 a_29161_n14476 0.020455f
C4881 a_27804_n14165 a_27700_n14116 0.026665f
C4882 a_27292_n14116 a_27496_n14116 0.048436f
C4883 a_42300_n13780 a_42188_n14213 0.026339f
C4884 a_23004_n2332 a_25975_n184 0.02831f
C4885 a_44092_n15348 VDD 0.3211f
C4886 a_47452_n2804 a_47900_n2804 0.012001f
C4887 a_22500_n1976 a_25084_1564 0.020992f
C4888 a_39164_n18484 VDD 0.319301f
C4889 a_24492_n5156 a_24180_n5112 0.464324f
C4890 a_41852_n4372 a_41740_n4805 0.026339f
C4891 a_34348_n17349 a_34796_n17349 0.012882f
C4892 a_41740_n6373 a_42188_n6373 0.012882f
C4893 a_30320_n6636 a_31936_n6592 0.011851f
C4894 a_47564_n7941 a_47476_n7844 0.285629f
C4895 a_38180_n20008 a_38628_n20008 0.013276f
C4896 a_45660_n2804 VDD 0.320877f
C4897 a_41292_n9509 a_41204_n9412 0.285629f
C4898 a_32132_2428 VDD 0.502437f
C4899 a_39500_n6373 VDD 0.319058f
C4900 a_39724_n11077 a_39636_n10980 0.285629f
C4901 a_46668_n9509 VDD 0.318039f
C4902 a_33488_n12996 a_34036_n12548 0.195478f
C4903 a_21772_n12996 a_21604_n13252 0.053827f
C4904 a_42636_n12645 a_43084_n12645 0.012882f
C4905 a_40396_n12645 VDD 0.334301f
C4906 a_21772_n12996 a_21604_n16872 0.017621f
C4907 a_40172_n15781 VDD 0.315469f
C4908 a_42188_n15781 a_42636_n15781 0.012882f
C4909 a_33900_n15781 a_33812_n15684 0.285629f
C4910 a_25084_1564 a_30296_1564 0.020914f
C4911 a_31324_n4372 a_31544_1248 0.059518f
C4912 a_30988_n18917 VDD 0.324804f
C4913 a_34796_n17349 a_35156_n17252 0.087066f
C4914 a_47116_n6373 a_47476_n6276 0.087066f
C4915 a_21604_n8548 a_22876_n8988 0.05539f
C4916 a_22016_n8961 a_22264_n8988 0.398421f
C4917 a_28335_n10644 a_27485_n10068 0.061094f
C4918 a_29532_n10311 a_29540_n11728 0.435107f
C4919 a_30604_1515 VDD 0.264767f
C4920 a_23016_n7376 VDD 0.36512f
C4921 a_47924_n4 VDD 0.213206f
C4922 a_42548_n10980 a_42996_n10980 0.013276f
C4923 a_26531_n10207 VDD 0.32564f
C4924 a_44876_n12645 a_44788_n12548 0.285629f
C4925 a_44788_n12548 VDD 0.22479f
C4926 a_40620_n14213 a_40532_n14116 0.285629f
C4927 a_32636_n2020 a_37632_n2020 0.181822f
C4928 a_44788_n15684 VDD 0.22479f
C4929 a_39948_n3237 a_40396_n3237 0.012001f
C4930 a_44428_n15781 a_44788_n15684 0.087066f
C4931 a_31544_1248 a_31961_1204 0.633318f
C4932 a_25972_n18820 VDD 0.209463f
C4933 a_28144_n4708 a_30215_n6265 0.033329f
C4934 a_45772_n17349 a_45684_n17252 0.285629f
C4935 a_40508_n4805 a_40420_n4708 0.285629f
C4936 a_35156_n17252 a_35604_n17252 0.013276f
C4937 a_23228_n6679 a_22772_n5808 0.027464f
C4938 a_22444_n5156 a_29612_n8292 0.023098f
C4939 a_45324_n101 VDD 0.323653f
C4940 a_24264_n6976 a_25685_n7463 0.015247f
C4941 a_23324_n7420 a_23220_n7376 0.026665f
C4942 a_30540_n18917 a_30452_n18820 0.285629f
C4943 a_22876_n4284 VDD 0.244849f
C4944 a_37844_n9412 a_37732_n10600 0.026657f
C4945 a_42212_n7464 VDD 0.206367f
C4946 a_24964_n14116 a_26239_n12996 0.045239f
C4947 a_26563_n12212 a_27055_n12168 0.092598f
C4948 a_42660_n18440 CLK 0.017841f
C4949 a_39972_n10600 VDD 0.207295f
C4950 a_46580_n12548 a_47028_n12548 0.013276f
C4951 a_45660_n1669 a_46108_n1669 0.013103f
C4952 a_31772_n16916 VDD 0.324283f
C4953 a_46580_n15684 a_47028_n15684 0.013276f
C4954 a_27337_n3140 a_28225_n4327 0.152423f
C4955 a_46668_n3237 a_47028_n3140 0.087066f
C4956 a_47476_n18820 VDD 0.206367f
C4957 a_41204_1243 a_42476_1515 0.05539f
C4958 a_45236_n4708 a_45684_n4708 0.013276f
C4959 a_41292_n18917 a_41652_n18820 0.087066f
C4960 a_33048_n7420 a_33497_n9032 0.047769f
C4961 a_27764_n18820 a_28212_n18820 0.013276f
C4962 a_42636_n9509 CLK 0.01698f
C4963 a_29444_n708 VDD 1.85667f
C4964 a_21604_n8548 a_23619_n9860 0.030097f
C4965 a_38180_n9032 a_38628_n9032 0.013276f
C4966 a_47116_n101 a_47564_n101 0.012222f
C4967 a_42660_n4328 VDD 0.206917f
C4968 a_25020_n11383 a_24964_n14116 0.038466f
C4969 a_30228_n8203 VDD 0.48537f
C4970 a_26547_n12951 VDD 0.604047f
C4971 a_43644_n13780 VDD 0.319164f
C4972 a_32308_n1976 a_34649_n2412 0.017545f
C4973 a_45572_n16872 VDD 0.213324f
C4974 a_22016_n4257 a_24128_n3840 0.277491f
C4975 a_23136_447 a_23728_464 0.869605f
C4976 a_33028_n20008 VDD 0.211234f
C4977 a_27092_n18440 a_27180_n18484 0.285629f
C4978 a_23036_n18484 a_23484_n18484 0.013103f
C4979 a_44004_n7464 a_44452_n7464 0.013276f
C4980 a_40420_n7464 a_40508_n7508 0.285629f
C4981 a_24672_n11339 a_25020_n11383 0.115314f
C4982 a_47364_n1192 VDD 0.206478f
C4983 a_25831_n11428 a_25237_n10599 0.090263f
C4984 a_28617_n8548 a_27281_n16854 0.023285f
C4985 a_37372_n20485 a_37732_n20388 0.087174f
C4986 a_25237_n5895 VDD 0.524996f
C4987 a_41764_n10600 a_42212_n10600 0.013276f
C4988 a_38180_n10600 a_38268_n10644 0.285629f
C4989 a_22220_n12996 a_22600_n12124 0.195081f
C4990 a_28437_n13705 a_24964_n14116 0.025076f
C4991 a_23564_n8292 a_23816_n13248 0.025372f
C4992 a_38068_n7844 VDD 0.230258f
C4993 a_45324_n11077 VDD 0.324845f
C4994 a_37859_377 a_41336_n407 0.028576f
C4995 a_35156_n13736 a_35604_n13736 0.013276f
C4996 a_22876_n1148 a_22568_n1104 0.934191f
C4997 a_22016_n1121 a_24233_n844 0.020455f
C4998 a_21604_n708 a_23816_n704 0.042802f
C4999 a_36140_n14213 VDD 0.296789f
C5000 a_26499_n2732 a_25895_n2624 0.387423f
C5001 a_35156_n15304 a_35244_n15348 0.285629f
C5002 a_27988_n4328 a_27932_n3543 0.022375f
C5003 a_43084_n17349 VDD 0.313885f
C5004 a_33564_n16916 a_34012_n16916 0.012552f
C5005 a_41864_1394 a_43101_841 0.018116f
C5006 a_39164_n20052 VDD 0.302205f
C5007 a_40980_n5896 a_41428_n5896 0.013276f
C5008 a_31236_n18440 a_30876_n18484 0.087066f
C5009 a_37732_n5896 a_37372_n5940 0.086742f
C5010 a_38180_n7464 CLK 0.0136f
C5011 a_46020_n7464 a_45660_n7508 0.086905f
C5012 a_29532_n10311 a_28435_n10599 0.017567f
C5013 a_44428_n4805 VDD 0.321554f
C5014 a_42748_n12212 a_43196_n12212 0.012882f
C5015 a_33910_n12146 a_34572_n12645 0.020327f
C5016 a_48012_332 a_48012_n101 0.05841f
C5017 a_39076_n13736 a_38716_n13780 0.087066f
C5018 a_29444_n708 a_31656_n704 0.042802f
C5019 a_30204_n1104 a_30408_n1104 0.048436f
C5020 a_46220_n101 a_46132_n4 0.285629f
C5021 a_40532_n14116 VDD 0.212412f
C5022 a_42660_n15304 a_43108_n15304 0.013276f
C5023 a_39076_n15304 a_39164_n15348 0.285629f
C5024 a_37221_n3543 a_35800_n3456 0.015898f
C5025 a_43892_n17252 VDD 0.210071f
C5026 a_40868_n16872 a_40508_n16916 0.087066f
C5027 a_40868_n4328 a_40508_n4372 0.087174f
C5028 a_23564_n20836 a_23484_n18484 0.013121f
C5029 a_34908_n20485 VDD 0.296789f
C5030 a_22588_n18484 a_22588_n18917 0.05841f
C5031 a_37732_n18440 a_38180_n18440 0.013276f
C5032 a_28324_n20008 a_27964_n20052 0.087066f
C5033 a_30228_n8203 a_30676_n7844 0.194599f
C5034 a_43780_n1572 VDD 0.20633f
C5035 a_26266_n9240 a_25724_n14564 0.022005f
C5036 a_24233_n5548 VDD 0.495722f
C5037 a_26547_n12951 a_27167_n10808 0.057143f
C5038 a_38716_n9076 VDD 0.321613f
C5039 a_28300_n15348 a_31664_n13292 0.037444f
C5040 a_21872_n12530 a_24573_n12996 0.463136f
C5041 a_37372_n12212 a_37260_n12645 0.026339f
C5042 a_38628_n12168 VDD 0.214363f
C5043 a_22600_n12124 a_23396_n16872 0.014067f
C5044 a_45572_n13736 a_46020_n13736 0.013276f
C5045 a_36052_n15304 VDD 0.203482f
C5046 a_27452_n2716 a_28583_n3140 0.27883f
C5047 a_43332_n2760 a_42972_n2804 0.087174f
C5048 a_27988_n4328 a_27540_n3797 0.20789f
C5049 a_27628_n3841 a_27932_n3543 0.039146f
C5050 a_32580_n18440 VDD 0.210284f
C5051 a_46020_n16872 a_46108_n16916 0.285629f
C5052 a_47364_n16872 a_47812_n16872 0.013276f
C5053 a_46020_n4328 a_45660_n4372 0.086905f
C5054 a_35268_n20388 VDD 0.203482f
C5055 a_39352_464 a_39804_464 0.026665f
C5056 a_25612_n6679 a_25524_n6635 0.494543f
C5057 a_29980_n18484 a_30092_n18917 0.026339f
C5058 a_31236_n20008 a_31324_n20052 0.285629f
C5059 a_34820_n20008 a_35268_n20008 0.013276f
C5060 a_36364_n7941 a_36276_n7844 0.285629f
C5061 a_33292_n2716 VDD 0.245641f
C5062 a_37484_n9509 a_37932_n9509 0.013103f
C5063 a_42860_n5940 VDD 0.329378f
C5064 a_30871_n11728 a_35716_n12168 0.020571f
C5065 a_46556_n12212 a_46668_n12645 0.026339f
C5066 a_42660_n20008 CLK 0.017841f
C5067 a_47812_n1192 a_47900_n1236 0.285629f
C5068 a_46108_n1236 a_46556_n1236 0.012552f
C5069 a_27804_n14165 a_27496_n14116 0.934191f
C5070 a_26944_n14116 a_28744_n14432 0.510371f
C5071 a_43644_n15348 VDD 0.319164f
C5072 a_44092_n15348 a_43980_n15781 0.026339f
C5073 a_38716_n18484 VDD 0.321613f
C5074 a_23887_n5156 a_24180_n5112 0.019052f
C5075 a_23207_n4708 a_23228_n6679 0.241041f
C5076 a_21692_n18917 a_22140_n18917 0.013103f
C5077 a_35916_n4 a_36120_n4 0.048436f
C5078 a_39860_n7844 a_40308_n7844 0.013276f
C5079 a_47116_n7941 a_47476_n7844 0.087066f
C5080 VDD OUT[5] 1.19171f
C5081 a_45212_n2804 VDD 0.343759f
C5082 a_40620_n9509 a_41204_n9412 0.016748f
C5083 a_47116_n11077 a_47564_n11077 0.012882f
C5084 a_39276_n11077 a_39636_n10980 0.087174f
C5085 a_46220_n9509 VDD 0.31977f
C5086 a_39948_n12645 VDD 0.31608f
C5087 a_37932_n14213 a_38380_n14213 0.012882f
C5088 a_39724_n15781 VDD 0.318714f
C5089 a_27628_n3841 a_27540_n3797 0.484626f
C5090 a_33452_n15781 a_33812_n15684 0.087066f
C5091 a_27988_n4328 a_27414_n5112 0.031544f
C5092 a_30540_n18917 VDD 0.321813f
C5093 a_34796_n17349 a_34708_n17252 0.285629f
C5094 a_44876_n17349 a_45324_n17349 0.012882f
C5095 a_41652_n6276 a_42100_n6276 0.013276f
C5096 a_46108_n18484 a_46220_n18917 0.026339f
C5097 a_47116_n6373 a_47028_n6276 0.285629f
C5098 a_25612_n6679 a_32856_n7376 0.029558f
C5099 a_42660_n9032 CLK 0.017841f
C5100 a_40956_n20052 a_41404_n20052 0.012882f
C5101 a_21604_n8548 a_22264_n8988 0.105778f
C5102 a_43892_n9412 a_44340_n9412 0.013276f
C5103 a_29992_n11150 a_30808_n10600 0.027343f
C5104 a_28836_376 VDD 0.614866f
C5105 a_22812_n7376 VDD 0.010384f
C5106 a_25412_n10600 VDD 0.124006f
C5107 a_35380_n12548 a_35828_n12548 0.013276f
C5108 a_44428_n12645 a_44788_n12548 0.087066f
C5109 a_44340_n12548 VDD 0.212126f
C5110 a_32308_n1572 a_32308_n1976 0.012806f
C5111 a_40172_n14213 a_40532_n14116 0.086635f
C5112 a_32636_n2020 a_36388_n1572 0.804001f
C5113 a_44340_n15684 VDD 0.212126f
C5114 a_44428_n15781 a_44340_n15684 0.285629f
C5115 a_35604_n15684 a_36052_n15684 0.013276f
C5116 a_25524_n18820 VDD 0.232671f
C5117 a_21692_2431 a_28132_376 0.033981f
C5118 a_45324_n17349 a_45684_n17252 0.087066f
C5119 a_40060_n4805 a_40420_n4708 0.086742f
C5120 a_46220_n4805 a_46668_n4805 0.012882f
C5121 a_42948_n1976 VDD 0.733446f
C5122 a_43532_n18917 a_43980_n18917 0.012882f
C5123 a_24681_n7116 a_25685_n7463 0.122205f
C5124 a_30092_n18917 a_30452_n18820 0.087066f
C5125 a_39164_n20052 a_39164_n20485 0.05841f
C5126 a_21792_n7464 VDD 0.505001f
C5127 a_26861_n10135 a_26239_n11428 0.022272f
C5128 a_25860_n9032 a_25880_n11708 0.487223f
C5129 a_41764_n7464 VDD 0.206367f
C5130 a_22904_n12080 a_23108_n12080 0.66083f
C5131 a_24964_n14116 a_25831_n12996 1.36977f
C5132 a_26563_n12212 a_26431_n12168 0.466019f
C5133 a_39524_n10600 VDD 0.209499f
C5134 a_42212_n18440 CLK 0.037136f
C5135 a_31455_n13648 VDD 0.046786f
C5136 a_42548_n14116 a_42996_n14116 0.013276f
C5137 a_32860_n2020 a_22820_n2804 0.193772f
C5138 a_31324_n4372 a_30716_n1148 0.013525f
C5139 a_31324_n16916 VDD 0.353532f
C5140 a_46668_n3237 a_46580_n3140 0.285629f
C5141 a_42100_n3140 a_42548_n3140 0.013276f
C5142 a_47028_n18820 VDD 0.206367f
C5143 a_41204_1243 a_41864_1394 0.108957f
C5144 a_45684_n17252 a_46132_n17252 0.013276f
C5145 a_23564_n20836 a_24380_n20052 0.012909f
C5146 a_29332_n17252 a_29444_n18440 0.026657f
C5147 a_41292_n18917 a_41204_n18820 0.285629f
C5148 a_24492_n5156 a_28868_n9387 0.011011f
C5149 a_23479_n5156 a_22220_n12996 0.027575f
C5150 a_32455_n7420 a_33497_n9032 0.354323f
C5151 a_42188_n9509 CLK 0.047331f
C5152 a_36924_n20485 a_37372_n20485 0.013103f
C5153 a_24604_n20485 a_24516_n20388 0.285629f
C5154 a_44509_n452 a_45236_n4 0.169257f
C5155 a_29532_n10311 a_22220_n12996 0.211172f
C5156 a_42212_n4328 VDD 0.206917f
C5157 a_28764_n8247 VDD 0.403145f
C5158 a_24964_n14116 VDD 0.998223f
C5159 a_38964_n12548 a_39076_n13736 0.026657f
C5160 a_43196_n13780 VDD 0.316157f
C5161 a_45572_n1572 a_46020_n1572 0.013276f
C5162 a_37396_n14116 a_37284_n15304 0.026657f
C5163 a_24220_n15260 a_25160_n14816 0.056721f
C5164 a_27192_n14286 a_27709_n16132 0.016134f
C5165 a_45124_n16872 VDD 0.26277f
C5166 a_40084_n15684 a_39972_n16872 0.026657f
C5167 a_32580_n20008 VDD 0.210015f
C5168 a_23136_447 a_24041_816 0.317251f
C5169 a_40420_n7464 a_40060_n7508 0.087066f
C5170 a_24292_n18820 a_24292_n20008 0.05841f
C5171 a_38292_n18820 a_38740_n18820 0.013276f
C5172 a_46916_n1192 VDD 0.206662f
C5173 a_40508_n9076 a_40956_n9076 0.012882f
C5174 a_37372_n20485 a_37284_n20388 0.285629f
C5175 a_24672_n11339 VDD 1.41986f
C5176 a_26239_n11428 a_26543_n11384 0.133465f
C5177 a_27281_n16854 a_26563_n12212 0.637858f
C5178 a_38180_n10600 a_37820_n10644 0.087066f
C5179 a_22220_n12996 a_22352_n12097 0.032445f
C5180 a_37620_n7844 VDD 0.213356f
C5181 a_40420_n12168 a_40868_n12168 0.013276f
C5182 a_44876_n11077 VDD 0.360805f
C5183 a_21604_n708 a_24233_n844 0.019043f
C5184 a_32152_n13692 a_33280_n13248 0.048436f
C5185 a_46132_n12548 a_46020_n13736 0.026657f
C5186 a_35692_n14213 VDD 0.296789f
C5187 a_25547_n2445 a_27348_n2672 0.427756f
C5188 a_32860_n2020 a_25237_n4327 1.48418f
C5189 a_35156_n15304 a_34796_n15348 0.087174f
C5190 a_42636_n17349 VDD 0.313885f
C5191 a_47028_n15684 a_46916_n16872 0.026657f
C5192 a_38716_n20052 VDD 0.304516f
C5193 a_41864_1394 a_42771_769 0.018275f
C5194 a_34372_n18440 a_34820_n18440 0.013276f
C5195 a_37284_n5896 a_37372_n5940 0.285629f
C5196 a_30788_n18440 a_30876_n18484 0.285629f
C5197 a_23564_n20836 a_24604_n20485 0.014129f
C5198 a_37732_n7464 CLK 0.0136f
C5199 a_46916_n7464 a_47364_n7464 0.013276f
C5200 a_31348_n18820 a_31236_n20008 0.026657f
C5201 a_24492_n5156 a_28927_n10160 0.019508f
C5202 a_45572_n7464 a_45660_n7508 0.285629f
C5203 a_37284_n20388 a_37732_n20388 0.013276f
C5204 a_25573_n12167 a_28335_n10644 0.036361f
C5205 a_25860_n9032 a_25020_n11383 0.041814f
C5206 a_43980_n4805 VDD 0.31896f
C5207 a_44540_n10644 a_45124_n10600 0.016748f
C5208 a_27281_n16854 a_27988_n20388 0.322741f
C5209 a_22904_n12080 VDD 0.364526f
C5210 a_30716_n1148 a_30408_n1104 0.934191f
C5211 a_42212_n13736 a_42660_n13736 0.013276f
C5212 a_38628_n13736 a_38716_n13780 0.285629f
C5213 a_29444_n708 a_32073_n844 0.019043f
C5214 a_45772_n101 a_46132_n4 0.086905f
C5215 a_40084_n14116 VDD 0.206509f
C5216 a_39076_n15304 a_38716_n15348 0.087066f
C5217 a_32432_n2689 a_34544_n2272 0.277491f
C5218 a_43444_n17252 VDD 0.208665f
C5219 a_25423_n4328 a_25530_n5112 0.016474f
C5220 a_40420_n4328 a_40508_n4372 0.285629f
C5221 a_40420_n16872 a_40508_n16916 0.285629f
C5222 a_44004_n16872 a_44452_n16872 0.013276f
C5223 a_34460_n20485 VDD 0.296789f
C5224 a_29612_n8292 a_29559_n6456 0.053278f
C5225 a_45124_n5896 a_45572_n5896 0.013276f
C5226 a_23564_n20836 a_24516_n20388 0.041882f
C5227 a_28764_n8247 a_30676_n7844 0.032459f
C5228 a_27876_n20008 a_27964_n20052 0.285629f
C5229 a_38292_n18820 a_38180_n20008 0.026657f
C5230 a_23932_n20052 a_24380_n20052 0.012882f
C5231 a_43332_n1572 VDD 0.196067f
C5232 a_25642_n9816 a_25724_n14564 0.021356f
C5233 a_25573_n12167 a_26239_n11428 0.021535f
C5234 a_44540_n9076 a_44428_n9509 0.026339f
C5235 a_40508_n10644 a_40620_n11077 0.026339f
C5236 a_38268_n9076 VDD 0.356786f
C5237 a_21872_n12530 a_23949_n12996 0.070346f
C5238 a_22600_n12124 a_22364_n13648 0.027048f
C5239 a_38180_n12168 VDD 0.245129f
C5240 a_22600_n12124 a_22948_n16872 0.015022f
C5241 a_34796_n13780 a_34796_n14213 0.05841f
C5242 a_35604_n15304 VDD 0.203482f
C5243 a_45572_n15304 a_46020_n15304 0.013276f
C5244 a_42884_n2760 a_42972_n2804 0.285629f
C5245 a_27988_n4328 a_28144_n4708 0.333134f
C5246 a_32132_n18440 VDD 0.212402f
C5247 a_46020_n16872 a_45660_n16916 0.086905f
C5248 a_45572_n4328 a_45660_n4372 0.285629f
C5249 a_46916_n4328 a_47364_n4328 0.013276f
C5250 a_24631_n3588 a_28548_n5112 0.032521f
C5251 a_34820_n20388 VDD 0.203482f
C5252 a_40508_n18484 a_40956_n18484 0.012882f
C5253 a_24573_n6724 a_25524_n6635 0.019347f
C5254 a_44452_n18440 a_44540_n18484 0.285629f
C5255 a_31236_n20008 a_30876_n20052 0.087066f
C5256 a_45236_n18820 a_45124_n20008 0.026657f
C5257 a_43084_n7941 a_43532_n7941 0.012882f
C5258 a_24492_n5156 a_29332_n11301 0.051874f
C5259 a_32432_n2689 VDD 0.800161f
C5260 a_42412_n5940 VDD 0.329378f
C5261 a_30871_n11728 a_35268_n12168 0.029678f
C5262 a_30428_n12645 a_30340_n12548 0.285629f
C5263 a_42212_n20008 CLK 0.037136f
C5264 a_47900_n12212 VDD 0.335152f
C5265 a_47812_n1192 a_47452_n1236 0.086635f
C5266 a_41852_n13780 a_41740_n14213 0.026339f
C5267 a_33252_n1192 a_33375_n1976 0.015261f
C5268 a_43196_n15348 VDD 0.316157f
C5269 a_47004_n2804 a_47452_n2804 0.012222f
C5270 a_38268_n18484 VDD 0.356784f
C5271 a_32132_2428 a_25084_1564 0.011005f
C5272 a_27988_n20388 a_27764_n18820 0.057406f
C5273 a_41404_n4372 a_41292_n4805 0.026339f
C5274 a_33900_n17349 a_34348_n17349 0.012882f
C5275 a_41292_n6373 a_41740_n6373 0.012882f
C5276 a_36428_n53 a_36120_n4 0.934191f
C5277 a_37732_n20008 a_38180_n20008 0.013276f
C5278 a_47116_n7941 a_47028_n7844 0.285629f
C5279 a_47116_n101 a_47028_n4 0.285629f
C5280 a_47812_n2760 VDD 0.209236f
C5281 a_40620_n9509 a_40532_n9412 0.285629f
C5282 a_22220_n12996 a_22568_n10512 0.015967f
C5283 a_25573_n12167 a_24684_n16432 0.38821f
C5284 a_30740_n7464 VDD 0.497292f
C5285 a_39276_n11077 a_39188_n10980 0.285629f
C5286 a_45772_n9509 VDD 0.321879f
C5287 a_42188_n12645 a_42636_n12645 0.012882f
C5288 a_39500_n12645 VDD 0.318341f
C5289 a_26271_n1400 a_26495_n1976 0.538085f
C5290 a_33077_n1191 a_34953_n1572 0.041737f
C5291 a_39276_n15781 VDD 0.320362f
C5292 a_41740_n15781 a_42188_n15781 0.012882f
C5293 a_27628_n3841 a_28144_n4708 0.16225f
C5294 a_33452_n15781 a_33364_n15684 0.285629f
C5295 a_25084_1564 a_30604_1515 0.018764f
C5296 a_30092_n18917 VDD 0.319783f
C5297 a_28548_n5112 a_30174_n5112 0.011071f
C5298 a_34348_n17349 a_34708_n17252 0.087066f
C5299 a_46668_n6373 a_47028_n6276 0.087066f
C5300 a_32332_n18917 a_32780_n18917 0.012001f
C5301 a_42212_n9032 CLK 0.037136f
C5302 a_21604_n8548 a_22016_n8961 0.536965f
C5303 a_29744_1564 VDD 0.824554f
C5304 a_23324_n7420 VDD 0.250021f
C5305 a_42100_n10980 a_42548_n10980 0.013276f
C5306 a_23816_n10112 VDD 1.37001f
C5307 a_44428_n12645 a_44340_n12548 0.285629f
C5308 a_43892_n12548 VDD 0.210071f
C5309 a_32636_n2020 a_36744_n1954 0.023664f
C5310 a_40172_n14213 a_40084_n14116 0.285629f
C5311 a_43892_n15684 VDD 0.210071f
C5312 a_43980_n15781 a_44340_n15684 0.087066f
C5313 a_39500_n3237 a_39948_n3237 0.012222f
C5314 a_21692_2431 a_28492_332 0.040641f
C5315 a_37859_377 a_40652_n1572 0.051291f
C5316 a_24740_n18820 VDD 0.241694f
C5317 a_45324_n17349 a_45236_n17252 0.285629f
C5318 a_40060_n4805 a_39972_n4708 0.285629f
C5319 a_34708_n17252 a_35156_n17252 0.013276f
C5320 a_22220_n9860 a_23816_n5408 0.038921f
C5321 a_44509_n452 VDD 0.735858f
C5322 a_37820_n5940 CLK 0.029648f
C5323 a_30092_n18917 a_30004_n18820 0.285629f
C5324 a_24681_n7116 a_24264_n6976 0.633318f
C5325 a_27485_n8500 a_28225_n9031 0.056162f
C5326 a_44340_n7844 a_44452_n9032 0.026657f
C5327 a_22016_n4257 VDD 0.804013f
C5328 a_37396_n9412 a_37284_n10600 0.026657f
C5329 a_45012_1564 VDD 0.164804f
C5330 a_26531_n10207 a_26239_n11428 0.216644f
C5331 a_41316_n7464 VDD 0.206367f
C5332 a_24684_n16432 a_21772_n12996 0.25617f
C5333 a_21772_n9860 a_27192_n14286 0.010001f
C5334 a_39076_n10600 VDD 0.211414f
C5335 a_46132_n12548 a_46580_n12548 0.013276f
C5336 a_32152_n13692 VDD 0.366412f
C5337 a_45212_n1669 a_45660_n1669 0.013103f
C5338 a_31324_n4372 a_29856_n1121 0.051284f
C5339 a_30876_n16916 VDD 0.323565f
C5340 a_27628_n3841 a_27190_n5112 0.010501f
C5341 a_46132_n15684 a_46580_n15684 0.013276f
C5342 a_46220_n3237 a_46580_n3140 0.087066f
C5343 a_41204_1243 a_41616_1564 0.536965f
C5344 a_46580_n18820 VDD 0.209166f
C5345 a_23564_n20836 a_23932_n20052 0.080406f
C5346 a_44788_n4708 a_45236_n4708 0.013276f
C5347 a_27316_n18820 a_27764_n18820 0.013276f
C5348 a_32560_n7020 a_33497_n9032 0.101226f
C5349 a_40620_n18917 a_41204_n18820 0.016748f
C5350 a_23479_n5156 a_26983_n12728 0.088378f
C5351 a_37732_n9032 a_38180_n9032 0.013276f
C5352 a_46668_n101 a_47116_n101 0.012222f
C5353 a_41764_n4328 VDD 0.206917f
C5354 a_32732_n10556 a_33672_n10112 0.056721f
C5355 a_25020_n11383 a_24760_n11383 0.484729f
C5356 a_28927_n10160 a_31664_n13292 0.01276f
C5357 a_42748_n13780 VDD 0.315469f
C5358 a_23608_n15260 a_25160_n14816 0.017769f
C5359 a_27192_n14286 a_27085_n16132 0.032639f
C5360 a_44540_n16916 VDD 0.353322f
C5361 a_32132_n20008 VDD 0.212133f
C5362 a_23136_447 a_23404_816 0.444933f
C5363 a_26084_n18440 a_26172_n18484 0.285629f
C5364 a_22588_n18484 a_23036_n18484 0.013103f
C5365 a_43556_n7464 a_44004_n7464 0.013276f
C5366 a_24492_n5156 a_25020_n11383 0.029971f
C5367 a_39972_n7464 a_40060_n7508 0.285629f
C5368 a_46468_n1192 VDD 0.209366f
C5369 a_44452_n9032 a_44540_n9076 0.285629f
C5370 a_36924_n20485 a_37284_n20388 0.087174f
C5371 a_26239_n11428 a_26547_n12951 0.073534f
C5372 a_22220_n12996 a_21940_n11684 0.07833f
C5373 a_41316_n10600 a_41764_n10600 0.013276f
C5374 a_42604_n2020 VDD 1.32713f
C5375 a_37732_n10600 a_37820_n10644 0.285629f
C5376 a_37172_n7844 VDD 0.211229f
C5377 a_44428_n11077 VDD 0.321554f
C5378 a_31559_n13692 a_33280_n13248 0.401636f
C5379 a_34708_n13736 a_35156_n13736 0.013276f
C5380 a_35244_n14213 VDD 0.296789f
C5381 a_34708_n15304 a_34796_n15348 0.285629f
C5382 a_22820_n2804 a_30555_n2729 0.205508f
C5383 a_42188_n17349 VDD 0.313885f
C5384 a_36612_n16872 a_36700_n16916 0.285629f
C5385 a_33116_n16916 a_33564_n16916 0.013103f
C5386 a_41864_1394 a_40776_770 0.076711f
C5387 a_38268_n20052 VDD 0.338723f
C5388 a_22220_n9860 a_23016_n7376 0.012195f
C5389 a_22444_n5156 a_30036_n7464 0.013014f
C5390 a_30788_n18440 a_30428_n18484 0.087066f
C5391 a_40532_n5896 a_40980_n5896 0.013276f
C5392 a_43555_n452 VDD 0.330497f
C5393 a_37284_n7464 CLK 0.0136f
C5394 a_25972_n6276 a_25831_n11428 0.181441f
C5395 a_45572_n7464 a_45212_n7508 0.086905f
C5396 a_24492_n5156 a_28437_n13705 0.039114f
C5397 a_33375_n1976 VDD 0.789578f
C5398 a_43532_n4805 VDD 0.317216f
C5399 a_25860_n9032 VDD 0.587856f
C5400 a_42300_n12212 a_42748_n12212 0.012882f
C5401 a_33686_n11592 a_34124_n12645 0.023919f
C5402 a_28121_n10980 a_27820_n16432 1.08846f
C5403 a_42548_n18820 CLK 0.029747f
C5404 a_22700_n12080 VDD 0.010384f
C5405 a_38628_n13736 a_38268_n13780 0.087066f
C5406 a_29856_n1121 a_30408_n1104 0.361958f
C5407 a_39636_n14116 VDD 0.209407f
C5408 a_42212_n15304 a_42660_n15304 0.013276f
C5409 a_38628_n15304 a_38716_n15348 0.285629f
C5410 a_47812_n1572 a_47812_n2760 0.05841f
C5411 a_31076_376 a_34895_n1192 0.05479f
C5412 a_42996_n17252 VDD 0.205948f
C5413 a_28144_n4708 a_22444_n5156 0.389064f
C5414 a_40420_n16872 a_40060_n16916 0.087066f
C5415 a_40420_n4328 a_40060_n4372 0.087174f
C5416 a_44004_n4328 a_44452_n4328 0.013276f
C5417 a_34012_n20485 VDD 0.296789f
C5418 a_31076_376 a_30104_n1148 0.540172f
C5419 a_29612_n8292 a_29211_n6724 0.046815f
C5420 a_22140_n18484 a_22140_n18917 0.05841f
C5421 a_37284_n18440 a_37732_n18440 0.013276f
C5422 a_27876_n20008 a_27516_n20052 0.087066f
C5423 a_28764_n8247 a_28972_n8247 0.489708f
C5424 a_25237_n10599 a_25724_n14564 0.476812f
C5425 a_25573_n12167 a_25500_n10644 0.04226f
C5426 a_33900_n11428 a_33364_n11384 0.407472f
C5427 a_26543_n11384 a_25559_n10980 0.056162f
C5428 a_37820_n9076 VDD 0.322978f
C5429 a_28300_n15348 a_30903_n13780 0.026969f
C5430 a_21872_n12530 a_22264_n13692 0.463958f
C5431 a_23619_n12996 a_23949_n12996 0.538085f
C5432 a_37732_n12168 VDD 0.213126f
C5433 a_22600_n12124 a_22500_n16872 0.01994f
C5434 a_45124_n13736 a_45572_n13736 0.013276f
C5435 a_35156_n15304 VDD 0.203482f
C5436 a_30555_n2729 a_25237_n4327 0.08262f
C5437 a_42884_n2760 a_42524_n2804 0.087174f
C5438 a_36588_n15348 a_36588_n15781 0.05841f
C5439 a_31684_n18440 VDD 0.218192f
C5440 a_46916_n16872 a_47364_n16872 0.013276f
C5441 a_45572_n4328 a_45212_n4372 0.086905f
C5442 a_45572_n16872 a_45660_n16916 0.285629f
C5443 a_34372_n20388 VDD 0.203482f
C5444 a_43725_908 a_44452_376 0.168987f
C5445 a_40776_770 a_40672_864 0.086548f
C5446 a_29532_n18484 a_29644_n18917 0.026339f
C5447 a_44452_n18440 a_44092_n18484 0.086635f
C5448 a_34372_n20008 a_34820_n20008 0.013276f
C5449 a_30788_n20008 a_30876_n20052 0.285629f
C5450 a_31392_n2760 VDD 0.227095f
C5451 a_37036_n9509 a_37484_n9509 0.013103f
C5452 a_41964_n5940 VDD 0.329378f
C5453 a_30871_n11728 a_33910_n12146 0.276523f
C5454 a_42324_n4 VDD 0.126246f
C5455 a_46108_n12212 a_46220_n12645 0.026339f
C5456 a_47452_n12212 VDD 0.313885f
C5457 a_47364_n1192 a_47452_n1236 0.285629f
C5458 a_26532_n14437 a_25636_n14520 0.015976f
C5459 a_27192_n14286 a_27292_n14116 0.087057f
C5460 a_26944_n14116 a_27496_n14116 0.361958f
C5461 a_45660_n1236 a_46108_n1236 0.012552f
C5462 a_42748_n15348 VDD 0.315469f
C5463 a_43644_n15348 a_43532_n15781 0.026339f
C5464 a_37820_n18484 VDD 0.322978f
C5465 a_27988_n20388 a_27316_n18820 0.014911f
C5466 a_27988_n4328 a_28121_n10980 0.055323f
C5467 a_46668_n7941 a_47028_n7844 0.087066f
C5468 a_39412_n7844 a_39860_n7844 0.013276f
C5469 a_46668_n101 a_47028_n4 0.086742f
C5470 a_47364_n2760 VDD 0.203482f
C5471 a_40172_n9509 a_40532_n9412 0.086742f
C5472 a_22220_n12996 a_22364_n10512 0.025643f
C5473 a_25573_n12167 a_25559_n10980 0.029138f
C5474 a_31068_n6276 VDD 0.31412f
C5475 a_46668_n11077 a_47116_n11077 0.012882f
C5476 a_24965_n9860 a_25642_n13736 0.032462f
C5477 a_38828_n11077 a_39188_n10980 0.087174f
C5478 a_45324_n9509 VDD 0.324845f
C5479 a_39052_n12645 VDD 0.320337f
C5480 a_37484_n14213 a_37932_n14213 0.012882f
C5481 a_38828_n15781 VDD 0.322604f
C5482 a_29644_n18917 VDD 0.317158f
C5483 a_25084_1564 a_28836_376 0.115718f
C5484 a_44428_n17349 a_44876_n17349 0.012882f
C5485 a_34348_n17349 a_34260_n17252 0.285629f
C5486 a_28548_n5112 a_29980_n5112 0.010472f
C5487 a_45660_n18484 a_45772_n18917 0.026339f
C5488 a_41204_n6276 a_41652_n6276 0.013276f
C5489 a_46668_n6373 a_46580_n6276 0.285629f
C5490 a_40508_n20052 a_40956_n20052 0.012882f
C5491 a_44452_n20008 a_44540_n20052 0.285629f
C5492 a_43444_n9412 a_43892_n9412 0.013276f
C5493 a_22712_n7420 VDD 0.731532f
C5494 a_24233_n10252 VDD 0.501519f
C5495 a_43980_n12645 a_44340_n12548 0.087066f
C5496 a_34932_n12548 a_35380_n12548 0.013276f
C5497 a_43444_n12548 VDD 0.208665f
C5498 a_39724_n14213 a_40084_n14116 0.087066f
C5499 a_32636_n2020 a_35940_n1931 0.013533f
C5500 a_43444_n15684 VDD 0.208665f
C5501 a_43980_n15781 a_43892_n15684 0.285629f
C5502 a_35156_n15684 a_35604_n15684 0.013276f
C5503 a_41864_1394 a_42772_n4 0.042966f
C5504 a_22500_n1976 a_23404_816 0.029217f
C5505 a_24292_n18820 VDD 0.212186f
C5506 a_39612_n4805 a_39972_n4708 0.086742f
C5507 a_45772_n4805 a_46220_n4805 0.012882f
C5508 a_22220_n9860 a_24233_n5548 0.0359f
C5509 a_44876_n17349 a_45236_n17252 0.087066f
C5510 a_28144_n4708 a_30320_n6636 0.022604f
C5511 a_43885_n452 VDD 0.583125f
C5512 a_37372_n5940 CLK 0.029648f
C5513 a_43084_n18917 a_43532_n18917 0.012882f
C5514 a_22464_n7393 a_24576_n6976 0.277491f
C5515 a_27988_n4328 a_29540_n11728 0.043075f
C5516 a_29644_n18917 a_30004_n18820 0.087066f
C5517 a_38716_n20052 a_38716_n20485 0.05841f
C5518 a_21604_n3844 VDD 1.81458f
C5519 a_43644_n705 VDD 1.35317f
C5520 a_40868_n7464 VDD 0.209318f
C5521 a_23212_n12124 a_23108_n12080 0.026665f
C5522 a_38628_n10600 VDD 0.214363f
C5523 a_31559_n13692 VDD 0.829307f
C5524 a_48012_n101 a_47924_n4 0.285629f
C5525 a_42100_n14116 a_42548_n14116 0.013276f
C5526 a_32132_2428 OUT[0] 0.022541f
C5527 a_30428_n16916 VDD 0.326298f
C5528 a_46220_n3237 a_46132_n3140 0.285629f
C5529 a_41652_n3140 a_42100_n3140 0.013276f
C5530 a_24631_n3588 a_25600_n5895 1.57746f
C5531 a_46132_n18820 VDD 0.210662f
C5532 a_45236_n17252 a_45684_n17252 0.013276f
C5533 a_23564_n20836 a_23484_n20052 0.043106f
C5534 a_40620_n18917 a_40532_n18820 0.285629f
C5535 a_33048_n7420 a_32856_n7376 0.934191f
C5536 a_35156_n325 a_35916_n4 0.011851f
C5537 a_23479_n5156 a_26635_n12996 0.071529f
C5538 a_41316_n4328 VDD 0.206917f
C5539 a_31872_n10529 a_33672_n10112 0.510371f
C5540 a_28435_n10599 a_33900_n11428 0.036237f
C5541 a_27597_n8292 VDD 0.733645f
C5542 a_24760_n11383 VDD 0.570102f
C5543 a_38516_n12548 a_38628_n13736 0.026657f
C5544 a_42300_n13780 VDD 0.315469f
C5545 a_23360_n15233 a_25160_n14816 0.510371f
C5546 a_45124_n1572 a_45572_n1572 0.013276f
C5547 a_44092_n16916 VDD 0.3211f
C5548 a_22876_n4284 a_23816_n3840 0.056721f
C5549 a_39636_n15684 a_39524_n16872 0.026657f
C5550 a_31684_n20008 VDD 0.217923f
C5551 a_26084_n18440 a_25724_n18484 0.086635f
C5552 a_23844_n18820 a_23844_n20008 0.05841f
C5553 a_37844_n18820 a_38292_n18820 0.013276f
C5554 a_39972_n7464 a_39612_n7508 0.087066f
C5555 a_46020_n1192 VDD 0.210709f
C5556 a_44452_n9032 a_44092_n9076 0.086635f
C5557 a_40060_n9076 a_40508_n9076 0.012882f
C5558 a_36924_n20485 a_36836_n20388 0.285629f
C5559 a_24492_n5156 VDD 1.2f
C5560 a_37732_n10600 a_37372_n10644 0.087066f
C5561 a_45660_332 VDD 0.32749f
C5562 a_36724_n7844 VDD 0.211674f
C5563 a_39972_n12168 a_40420_n12168 0.013276f
C5564 a_43980_n11077 VDD 0.31896f
C5565 a_45684_n12548 a_45572_n13736 0.026657f
C5566 a_22016_n1121 a_22568_n1104 0.361958f
C5567 a_31664_n13292 a_33280_n13248 0.011851f
C5568 a_34796_n14213 VDD 0.296789f
C5569 a_34708_n15304 a_34348_n15348 0.087174f
C5570 a_23004_n2332 a_22568_n1104 0.031141f
C5571 a_41740_n17349 VDD 0.313885f
C5572 a_36612_n16872 a_36252_n16916 0.086635f
C5573 a_46580_n15684 a_46468_n16872 0.026657f
C5574 a_22052_n4708 a_23228_n6679 0.0272f
C5575 a_37820_n20052 VDD 0.305881f
C5576 a_30340_n18440 a_30428_n18484 0.285629f
C5577 a_22444_n5156 a_30396_n7508 0.019315f
C5578 a_33924_n18440 a_34372_n18440 0.013276f
C5579 a_42860_n101 VDD 0.333185f
C5580 a_30900_n18820 a_30788_n20008 0.026657f
C5581 a_46468_n7464 a_46916_n7464 0.013276f
C5582 a_25972_n6276 a_34092_n9076 0.241702f
C5583 a_45124_n7464 a_45212_n7508 0.285629f
C5584 a_32860_n2020 VDD 0.867248f
C5585 a_29532_n10311 a_28927_n10160 0.722238f
C5586 a_36836_n20388 a_37284_n20388 0.013276f
C5587 a_43084_n4805 VDD 0.313885f
C5588 a_44092_n10644 a_44540_n10644 0.012001f
C5589 a_25412_n8501 VDD 0.442403f
C5590 a_23212_n12124 VDD 0.248562f
C5591 a_42100_n18820 CLK 0.020589f
C5592 a_38180_n13736 a_38268_n13780 0.285629f
C5593 a_41764_n13736 a_42212_n13736 0.013276f
C5594 a_29856_n1121 a_30204_n1104 0.401636f
C5595 a_39188_n14116 VDD 0.211136f
C5596 a_38628_n15304 a_38268_n15348 0.087066f
C5597 a_31076_376 a_34271_n1192 0.46464f
C5598 a_42548_n17252 VDD 0.205948f
C5599 a_39972_n16872 a_40060_n16916 0.285629f
C5600 a_43556_n16872 a_44004_n16872 0.013276f
C5601 a_39972_n4328 a_40060_n4372 0.285629f
C5602 a_33564_n20485 VDD 0.296789f
C5603 a_27428_n20008 a_27516_n20052 0.285629f
C5604 a_37844_n18820 a_37732_n20008 0.026657f
C5605 a_23484_n20052 a_23932_n20052 0.012882f
C5606 a_44092_n9076 a_43980_n9509 0.026339f
C5607 a_24965_n9860 a_25724_n14564 0.659613f
C5608 a_22568_n5808 VDD 0.362268f
C5609 a_24964_n14116 a_24684_n16432 0.352667f
C5610 a_40060_n10644 a_40172_n11077 0.026339f
C5611 a_37372_n9076 VDD 0.327457f
C5612 a_21872_n12530 a_22116_n12548 0.014831f
C5613 a_23619_n12996 a_22264_n13692 0.234246f
C5614 a_22600_n12124 a_22016_n13665 0.047079f
C5615 a_37284_n12168 VDD 0.231657f
C5616 a_42157_n660 a_42884_n1192 0.168987f
C5617 a_34708_n15304 VDD 0.203482f
C5618 a_45124_n15304 a_45572_n15304 0.013276f
C5619 a_27452_n2716 a_25600_n5895 0.374063f
C5620 a_42436_n2760 a_42524_n2804 0.285629f
C5621 a_31236_n18440 VDD 0.22735f
C5622 a_45572_n16872 a_45212_n16916 0.086905f
C5623 a_46468_n4328 a_46916_n4328 0.013276f
C5624 a_45124_n4328 a_45212_n4372 0.285629f
C5625 a_39544_420 a_39804_464 0.66083f
C5626 a_43725_908 a_40260_n408 0.473675f
C5627 a_33924_n20388 VDD 0.203482f
C5628 a_44004_n18440 a_44092_n18484 0.285629f
C5629 a_40060_n18484 a_40508_n18484 0.012882f
C5630 a_42636_n7941 a_43084_n7941 0.012882f
C5631 a_31965_n8292 a_29532_n10311 0.12552f
C5632 a_30788_n20008 a_30428_n20052 0.087066f
C5633 a_31412_n2276 VDD 0.810335f
C5634 a_29532_n10311 a_29332_n11301 0.031097f
C5635 a_41516_n5940 VDD 0.329378f
C5636 a_35064_n11383 a_34350_n10980 0.484512f
C5637 a_30871_n11728 a_33686_n11592 0.043697f
C5638 a_28121_n10980 a_28752_n15348 0.02811f
C5639 a_47004_n12212 VDD 0.313885f
C5640 a_41404_n13780 a_41292_n14213 0.026339f
C5641 a_47364_n1192 a_47004_n1236 0.086742f
C5642 a_26944_n14116 a_27292_n14116 0.401636f
C5643 a_28132_376 a_26736_n364 0.036238f
C5644 a_42300_n15348 VDD 0.315469f
C5645 a_46556_n2804 a_47004_n2804 0.012222f
C5646 a_32132_2428 a_31324_n4372 0.585164f
C5647 a_22500_n1976 a_28736_1944 1.45455f
C5648 a_37372_n18484 VDD 0.324575f
C5649 a_33452_n17349 a_33900_n17349 0.012882f
C5650 a_24672_n11339 a_22220_n9860 1.39486f
C5651 a_46668_n7941 a_46580_n7844 0.285629f
C5652 a_37284_n20008 a_37732_n20008 0.013276f
C5653 a_46916_n2760 VDD 0.203495f
C5654 a_40172_n9509 a_40084_n9412 0.285629f
C5655 a_22220_n12996 a_22876_n10556 0.016287f
C5656 a_47564_n9509 a_48012_n9509 0.012882f
C5657 a_30616_n6221 VDD 0.261269f
C5658 a_26543_n11384 a_26431_n12168 0.026175f
C5659 a_24965_n9860 a_25237_n13735 0.046017f
C5660 a_38828_n11077 a_38740_n10980 0.285629f
C5661 a_44876_n9509 VDD 0.360805f
C5662 a_41740_n12645 a_42188_n12645 0.012882f
C5663 a_38604_n12645 VDD 0.322952f
C5664 a_38380_n15781 VDD 0.342527f
C5665 a_41292_n15781 a_41740_n15781 0.012882f
C5666 a_25084_1564 a_29744_1564 0.028467f
C5667 a_29196_n18917 VDD 0.330964f
C5668 a_33900_n17349 a_34260_n17252 0.087066f
C5669 a_31884_n18917 a_32332_n18917 0.012882f
C5670 a_46220_n6373 a_46580_n6276 0.087066f
C5671 a_25612_n6679 a_33048_n7420 0.016277f
C5672 a_44452_n20008 a_44092_n20052 0.086635f
C5673 a_22464_n7393 VDD 0.8193f
C5674 a_41652_n10980 a_42100_n10980 0.013276f
C5675 a_43980_n12645 a_43892_n12548 0.285629f
C5676 a_42996_n12548 VDD 0.205948f
C5677 a_39724_n14213 a_39636_n14116 0.285629f
C5678 a_33375_n1976 a_33999_n1400 0.104193f
C5679 a_42996_n15684 VDD 0.205948f
C5680 a_43532_n15781 a_43892_n15684 0.087066f
C5681 a_44004_n1192 a_41616_1564 0.012798f
C5682 a_23844_n18820 VDD 0.208184f
C5683 a_30296_1564 a_30500_1564 0.66083f
C5684 a_34260_n17252 a_34708_n17252 0.013276f
C5685 a_39612_n4805 a_39524_n4708 0.285629f
C5686 a_28144_n4708 a_29559_n6456 0.033963f
C5687 a_44876_n17349 a_44788_n17252 0.285629f
C5688 a_29644_n18917 a_29556_n18820 0.285629f
C5689 a_27988_n4328 a_28009_n12168 0.19616f
C5690 a_23564_n8292 a_22220_n12996 0.03094f
C5691 a_25573_n12167 a_28617_n8548 0.111403f
C5692 a_43892_n7844 a_44004_n9032 0.026657f
C5693 a_25412_n10600 a_25500_n10644 0.285629f
C5694 a_40420_n7464 VDD 0.206367f
C5695 a_24964_n14116 a_24573_n12996 0.039826f
C5696 a_38180_n10600 VDD 0.245129f
C5697 a_36120_n4 a_36324_n4 0.66083f
C5698 a_45684_n12548 a_46132_n12548 0.013276f
C5699 a_31664_n13292 VDD 1.80482f
C5700 a_47564_n101 a_47924_n4 0.086635f
C5701 VDD EOC 1.03725f
C5702 a_44764_n1669 a_45212_n1669 0.013103f
C5703 a_27988_n4328 a_22164_n2760 0.023816f
C5704 a_31324_n4372 a_29444_n708 0.015771f
C5705 a_36612_n16872 VDD 0.215878f
C5706 a_45772_n3237 a_46132_n3140 0.087066f
C5707 a_45684_n15684 a_46132_n15684 0.013276f
C5708 a_27932_n3543 a_28225_n4327 0.304801f
C5709 a_45684_n18820 VDD 0.212897f
C5710 a_44340_n4708 a_44788_n4708 0.013276f
C5711 a_40172_n18917 a_40532_n18820 0.086635f
C5712 a_26868_n18820 a_27316_n18820 0.013276f
C5713 a_32455_n7420 a_32856_n7376 0.882105f
C5714 a_35156_n325 a_36428_n53 0.05539f
C5715 a_37284_n9032 a_37732_n9032 0.013276f
C5716 a_23479_n5156 a_26239_n12996 0.033745f
C5717 a_46220_n101 a_46668_n101 0.012552f
C5718 a_40868_n4328 VDD 0.209985f
C5719 a_31872_n10529 a_34089_n10252 0.020455f
C5720 a_26973_n8292 VDD 0.581617f
C5721 a_25724_n14564 a_25636_n14520 0.521468f
C5722 a_28927_n10160 a_30903_n13780 0.016109f
C5723 a_23564_n11428 VDD 1.21515f
C5724 a_26563_n12212 a_27524_n15304 0.01472f
C5725 a_41852_n13780 VDD 0.315469f
C5726 a_23360_n15233 a_25577_n14956 0.020455f
C5727 a_23708_n15216 a_23912_n15216 0.048436f
C5728 a_43644_n16916 VDD 0.319164f
C5729 a_31236_n20008 VDD 0.226508f
C5730 a_27988_n4328 a_22220_n12996 0.037114f
C5731 a_22140_n18484 a_22588_n18484 0.013103f
C5732 a_25636_n18440 a_25724_n18484 0.285629f
C5733 a_39524_n7464 a_39612_n7508 0.285629f
C5734 a_23479_n5156 a_25020_n11383 0.043744f
C5735 a_26943_n7442 a_27597_n8292 0.017184f
C5736 a_43108_n7464 a_43556_n7464 0.013276f
C5737 a_45572_n1192 VDD 0.211391f
C5738 a_36252_n20485 a_36836_n20388 0.016748f
C5739 a_29532_n10311 a_25020_n11383 0.030791f
C5740 a_44004_n9032 a_44092_n9076 0.285629f
C5741 a_47228_n20485 a_47676_n20485 0.013103f
C5742 a_23887_n5156 VDD 0.733913f
C5743 a_25500_n10644 a_24964_n14116 0.018289f
C5744 a_37284_n10600 a_37372_n10644 0.285629f
C5745 a_40868_n10600 a_41316_n10600 0.013276f
C5746 a_45212_332 VDD 0.341634f
C5747 a_36276_n7844 VDD 0.145712f
C5748 a_43532_n11077 VDD 0.317216f
C5749 a_21604_n708 a_22568_n1104 0.08126f
C5750 a_22016_n1121 a_22364_n1104 0.401636f
C5751 a_34348_n14213 VDD 0.328124f
C5752 a_22164_n2760 a_27628_n3841 0.585126f
C5753 a_34260_n15304 a_34348_n15348 0.285629f
C5754 a_41292_n17349 VDD 0.318502f
C5755 a_32668_n16916 a_33116_n16916 0.013103f
C5756 a_36164_n16872 a_36252_n16916 0.285629f
C5757 a_37372_n20052 VDD 0.307479f
C5758 a_24492_n5156 a_26943_n7442 0.028017f
C5759 a_22220_n9860 a_23324_n7420 0.015841f
C5760 a_30340_n18440 a_29980_n18484 0.087066f
C5761 a_40084_n5896 a_40532_n5896 0.013276f
C5762 a_42412_n101 VDD 0.331075f
C5763 a_25972_n6276 a_33832_n8572 0.023868f
C5764 a_32636_n2020 VDD 0.448278f
C5765 a_47452_n9076 a_47900_n9076 0.012001f
C5766 a_47676_n20485 a_47588_n20388 0.285629f
C5767 a_42636_n4805 VDD 0.313885f
C5768 a_45236_n4 a_45124_n1192 0.026657f
C5769 a_22772_n8944 VDD 0.299247f
C5770 a_32854_n12168 a_33488_n12996 0.012015f
C5771 a_41852_n12212 a_42300_n12212 0.012882f
C5772 a_22600_n12124 VDD 0.73171f
C5773 a_38180_n13736 a_37820_n13780 0.087066f
C5774 a_29444_n708 a_30408_n1104 0.08126f
C5775 a_29856_n1121 a_30716_n1148 0.882105f
C5776 a_38740_n14116 VDD 0.213797f
C5777 a_38180_n15304 a_38268_n15348 0.285629f
C5778 a_33292_n2716 a_34232_n2272 0.056721f
C5779 a_47364_n1572 a_47364_n2760 0.05841f
C5780 a_41764_n15304 a_42212_n15304 0.013276f
C5781 a_42100_n17252 VDD 0.205948f
C5782 a_43556_n4328 a_44004_n4328 0.013276f
C5783 a_39972_n4328 a_39612_n4372 0.087174f
C5784 a_39972_n16872 a_39612_n16916 0.087066f
C5785 a_33116_n20485 VDD 0.303438f
C5786 a_21692_n18484 a_21692_n18917 0.05841f
C5787 a_36700_n18484 a_37284_n18440 0.016748f
C5788 a_28764_n8247 a_29176_n7819 0.025326f
C5789 a_27428_n20008 a_27068_n20052 0.087066f
C5790 a_44540_n7508 a_44428_n7941 0.026339f
C5791 a_41204_n1572 VDD 0.227989f
C5792 a_25860_n9032 a_26239_n11428 0.097306f
C5793 a_22364_n5808 VDD 0.010384f
C5794 a_24964_n14116 a_25559_n10980 0.077464f
C5795 a_24965_n9860 a_25132_n16432 0.315594f
C5796 a_28300_n15348 a_27820_n16432 0.023101f
C5797 a_36700_n12212 VDD 0.345602f
C5798 a_44540_n13780 a_45124_n13736 0.016748f
C5799 a_34260_n15304 VDD 0.203482f
C5800 a_36140_n15348 a_36140_n15781 0.05841f
C5801 a_42436_n2760 a_42076_n2804 0.087174f
C5802 a_30788_n18440 VDD 0.212672f
C5803 a_46468_n16872 a_46916_n16872 0.013276f
C5804 a_45124_n16872 a_45212_n16916 0.285629f
C5805 a_43101_841 a_40260_n408 0.093491f
C5806 a_33476_n20388 VDD 0.203482f
C5807 a_23949_n6724 a_24573_n6724 0.104193f
C5808 a_44004_n18440 a_43644_n18484 0.087066f
C5809 a_30340_n20008 a_30428_n20052 0.285629f
C5810 a_33924_n20008 a_34372_n20008 0.013276f
C5811 a_23479_n5156 a_27391_n11384 0.064949f
C5812 a_30555_n2729 VDD 1.01918f
C5813 a_36588_n9509 a_37036_n9509 0.013103f
C5814 a_41068_n5940 VDD 0.328713f
C5815 a_30871_n11728 a_32854_n12168 0.044348f
C5816 a_45660_n12212 a_45772_n12645 0.026339f
C5817 a_46556_n12212 VDD 0.31705f
C5818 a_26532_n14437 a_29161_n14476 0.019043f
C5819 a_26944_n14116 a_27804_n14165 0.882105f
C5820 a_46916_n1192 a_47004_n1236 0.285629f
C5821 a_45212_n1236 a_45660_n1236 0.012552f
C5822 a_31656_n704 a_32636_n2020 0.029124f
C5823 a_28492_332 a_26736_n364 0.030312f
C5824 a_41852_n15348 VDD 0.315469f
C5825 a_43196_n15348 a_43084_n15781 0.026339f
C5826 a_22500_n15684 a_22948_n15684 0.013276f
C5827 a_44452_n18440 VDD 0.219497f
C5828 a_40508_n4372 a_40508_n4805 0.05841f
C5829 a_26154_n4536 a_26358_n4618 0.499501f
C5830 a_47452_n18484 a_47900_n18484 0.012001f
C5831 a_42604_n2020 a_46132_n4 0.047963f
C5832 a_38964_n7844 a_39412_n7844 0.013276f
C5833 a_46220_n7941 a_46580_n7844 0.087066f
C5834 a_46468_n2760 VDD 0.206589f
C5835 a_22220_n12996 a_22016_n10529 0.081298f
C5836 a_39724_n9509 a_40084_n9412 0.086742f
C5837 a_25860_n9032 a_24684_n16432 0.010668f
C5838 a_26607_1966 VDD 0.309232f
C5839 a_30111_n6221 VDD 0.022335f
C5840 a_26547_n12951 a_26431_n12168 0.074818f
C5841 a_46220_n11077 a_46668_n11077 0.012882f
C5842 a_24965_n9860 a_23816_n13248 0.049678f
C5843 a_38380_n11077 a_38740_n10980 0.087174f
C5844 a_44428_n9509 VDD 0.321554f
C5845 a_38156_n12645 VDD 0.356085f
C5846 a_37036_n14213 a_37484_n14213 0.012882f
C5847 a_37932_n15781 VDD 0.327654f
C5848 a_28568_n16066 a_23564_n17700 0.432794f
C5849 a_44316_n2804 a_44428_n3237 0.026339f
C5850 a_32132_2428 a_31544_1248 0.022039f
C5851 a_28748_n18917 VDD 0.329708f
C5852 a_33900_n17349 a_33812_n17252 0.285629f
C5853 a_43980_n17349 a_44428_n17349 0.012882f
C5854 a_46220_n6373 a_46132_n6276 0.285629f
C5855 a_25612_n6679 a_32455_n7420 0.038517f
C5856 a_45212_n18484 a_45324_n18917 0.026339f
C5857 a_44004_n20008 a_44092_n20052 0.285629f
C5858 a_40060_n20052 a_40508_n20052 0.012882f
C5859 a_29532_n10311 a_32767_n9010 0.083656f
C5860 a_42996_n9412 a_43444_n9412 0.013276f
C5861 a_29332_1243 VDD 1.75962f
C5862 a_22052_n6980 VDD 1.75201f
C5863 a_43532_n12645 a_43892_n12548 0.087066f
C5864 a_34484_n12548 a_34932_n12548 0.013276f
C5865 a_42548_n12548 VDD 0.205948f
C5866 a_26532_n14437 a_27404_n14990 0.035919f
C5867 a_39276_n14213 a_39636_n14116 0.087066f
C5868 a_32636_n2020 a_34223_n1976 0.019338f
C5869 a_42548_n15684 VDD 0.205948f
C5870 a_34708_n15684 a_35156_n15684 0.013276f
C5871 a_43532_n15781 a_43444_n15684 0.285629f
C5872 a_29744_1564 a_31856_1248 0.277491f
C5873 a_30604_1515 a_31544_1248 0.056721f
C5874 a_23396_n18820 VDD 0.207289f
C5875 a_44428_n17349 a_44788_n17252 0.087066f
C5876 a_39164_n4805 a_39524_n4708 0.086905f
C5877 a_28144_n4708 a_29211_n6724 0.0132f
C5878 a_45324_n4805 a_45772_n4805 0.012882f
C5879 a_29196_n18917 a_29556_n18820 0.087066f
C5880 a_42636_n18917 a_43084_n18917 0.012882f
C5881 a_38268_n20052 a_38268_n20485 0.05841f
C5882 a_39972_n7464 VDD 0.207713f
C5883 a_24569_n11820 a_24152_n11680 0.633318f
C5884 a_37732_n10600 VDD 0.213126f
C5885 a_36428_n53 a_37368_n320 0.056721f
C5886 a_41652_n14116 a_42100_n14116 0.013276f
C5887 a_36164_n16872 VDD 0.207033f
C5888 a_45772_n3237 a_45684_n3140 0.285629f
C5889 a_41204_n3140 a_41652_n3140 0.013276f
C5890 a_24631_n3588 a_27337_n3140 0.039224f
C5891 a_45236_n18820 VDD 0.229931f
C5892 a_44788_n17252 a_45236_n17252 0.013276f
C5893 a_40172_n18917 a_40084_n18820 0.285629f
C5894 a_32560_n7020 a_32856_n7376 0.05539f
C5895 a_25524_n708 VDD 0.797281f
C5896 a_35804_n20485 a_36252_n20485 0.013103f
C5897 a_23479_n5156 a_25831_n12996 0.025532f
C5898 a_40420_n4328 VDD 0.206917f
C5899 a_28435_n10599 a_32628_n10512 0.014595f
C5900 a_32220_n10512 a_32424_n10512 0.048436f
C5901 a_31076_376 VDD 0.939952f
C5902 a_25132_n16432 a_25636_n14520 0.025079f
C5903 a_38068_n12548 a_38180_n13736 0.026657f
C5904 a_41404_n13780 VDD 0.315469f
C5905 a_44676_n1572 a_45124_n1572 0.013276f
C5906 a_24220_n15260 a_23912_n15216 0.934191f
C5907 a_43196_n16916 VDD 0.316157f
C5908 a_39188_n15684 a_39076_n16872 0.026657f
C5909 a_22016_n4257 a_23816_n3840 0.510371f
C5910 a_30788_n20008 VDD 0.212403f
C5911 a_25636_n18440 a_25276_n18484 0.086742f
C5912 a_23816_n5408 a_24128_n5408 0.119687f
C5913 a_24492_n5156 a_28335_n10644 0.026219f
C5914 a_23396_n18820 a_23396_n20008 0.05841f
C5915 a_39524_n7464 a_39164_n7508 0.087066f
C5916 a_37396_n18820 a_37844_n18820 0.013276f
C5917 a_45124_n1192 VDD 0.263858f
C5918 a_44004_n9032 a_43644_n9076 0.087066f
C5919 a_39612_n9076 a_40060_n9076 0.012882f
C5920 a_36252_n20485 a_36164_n20388 0.285629f
C5921 a_23479_n5156 VDD 1.38892f
C5922 a_47924_376 VDD 0.129633f
C5923 a_29532_n10311 VDD 1.1889f
C5924 a_39524_n12168 a_39972_n12168 0.013276f
C5925 a_43084_n11077 VDD 0.313885f
C5926 a_22016_n1121 a_22876_n1148 0.882105f
C5927 a_45236_n12548 a_45124_n13736 0.026657f
C5928 a_21604_n708 a_22364_n1104 0.011851f
C5929 a_33900_n14213 VDD 0.321896f
C5930 a_25547_n2445 a_27452_n2716 0.41094f
C5931 a_34260_n15304 a_33900_n15348 0.087174f
C5932 a_23004_n2332 a_22876_n1148 0.028326f
C5933 a_40620_n17349 VDD 0.343849f
C5934 a_46132_n15684 a_46020_n16872 0.026657f
C5935 a_28144_n4708 a_28225_n4327 0.052766f
C5936 a_36164_n16872 a_35804_n16916 0.086742f
C5937 a_22052_n4708 a_26358_n4618 0.014835f
C5938 a_44452_n20008 VDD 0.219497f
C5939 a_28492_332 a_32909_841 0.015207f
C5940 a_22220_n9860 a_22712_n7420 0.034478f
C5941 a_24492_n5156 a_26719_n7464 0.013469f
C5942 a_29892_n18440 a_29980_n18484 0.285629f
C5943 a_33476_n18440 a_33924_n18440 0.013276f
C5944 a_41336_n407 VDD 0.470388f
C5945 a_46020_n7464 a_46468_n7464 0.013276f
C5946 a_30452_n18820 a_30340_n20008 0.026657f
C5947 a_47228_n20485 a_47588_n20388 0.087174f
C5948 a_42188_n4805 VDD 0.313885f
C5949 a_43644_n10644 a_44092_n10644 0.012882f
C5950 a_24128_n8544 VDD 0.02612f
C5951 a_22352_n12097 VDD 0.809227f
C5952 a_37732_n13736 a_37820_n13780 0.285629f
C5953 a_41316_n13736 a_41764_n13736 0.013276f
C5954 a_29444_n708 a_30204_n1104 0.011851f
C5955 a_38292_n14116 VDD 0.243749f
C5956 a_38180_n15304 a_37820_n15348 0.087066f
C5957 a_32432_n2689 a_34232_n2272 0.510371f
C5958 a_41652_n17252 VDD 0.205948f
C5959 a_43108_n16872 a_43556_n16872 0.013276f
C5960 a_39524_n16872 a_39612_n16916 0.285629f
C5961 a_39524_n4328 a_39612_n4372 0.285629f
C5962 a_32444_n20485 VDD 0.362778f
C5963 a_43756_n5940 a_44204_n5940 0.012222f
C5964 a_26980_n20008 a_27068_n20052 0.285629f
C5965 a_37396_n18820 a_37284_n20008 0.026657f
C5966 a_23036_n20052 a_23484_n20052 0.012882f
C5967 a_43644_n9076 a_43532_n9509 0.026339f
C5968 a_22876_n5852 VDD 0.245825f
C5969 a_39612_n10644 a_39724_n11077 0.026339f
C5970 a_34652_n11391 a_28300_n15348 0.099078f
C5971 a_35119_398 a_35156_n325 0.030073f
C5972 a_44452_n9032 VDD 0.219497f
C5973 a_23619_n12996 a_21872_n12530 0.018938f
C5974 a_36252_n12212 VDD 0.313975f
C5975 a_41533_n727 a_42157_n660 0.104193f
C5976 a_33812_n15304 VDD 0.203482f
C5977 a_41988_n2760 a_42076_n2804 0.285629f
C5978 a_44540_n15348 a_45124_n15304 0.016748f
C5979 a_30340_n18440 VDD 0.210564f
C5980 a_46020_n4328 a_46468_n4328 0.013276f
C5981 a_43101_841 a_43725_908 0.104193f
C5982 a_33028_n20388 VDD 0.22685f
C5983 a_42771_769 a_40260_n408 0.031586f
C5984 a_43556_n18440 a_43644_n18484 0.285629f
C5985 a_39612_n18484 a_40060_n18484 0.012882f
C5986 a_23479_n5156 a_27167_n10808 0.06034f
C5987 a_30676_n7844 a_29532_n10311 0.020891f
C5988 a_42188_n7941 a_42636_n7941 0.012882f
C5989 a_30340_n20008 a_29980_n20052 0.087066f
C5990 a_40620_n5940 VDD 0.329378f
C5991 a_30871_n11728 a_32650_n12168 0.034809f
C5992 a_21892_n9816 VDD 0.824292f
C5993 a_46108_n12212 VDD 0.318654f
C5994 a_26532_n14437 a_28744_n14432 0.042802f
C5995 a_26944_n14116 a_27192_n14286 0.33448f
C5996 a_46916_n1192 a_46556_n1236 0.086742f
C5997 a_27572_860 a_26736_n364 0.035903f
C5998 a_41404_n15348 VDD 0.315469f
C5999 a_26755_n16132 a_27085_n16132 0.538085f
C6000 a_46108_n2804 a_46556_n2804 0.012552f
C6001 a_47812_n2760 a_47900_n2804 0.285629f
C6002 a_44004_n18440 VDD 0.2108f
C6003 a_24492_n5156 a_22220_n9860 0.156221f
C6004 a_22788_n4708 a_22564_n5112 0.013419f
C6005 a_46132_n4 a_46020_n1192 0.026657f
C6006 a_39948_n6373 a_40396_n6373 0.012001f
C6007 a_36700_n20052 a_37284_n20008 0.016748f
C6008 a_46220_n7941 a_46132_n7844 0.285629f
C6009 a_46020_n2760 VDD 0.20827f
C6010 a_39724_n9509 a_39636_n9412 0.285629f
C6011 a_22220_n12996 a_21604_n10116 0.011407f
C6012 a_47116_n9509 a_47564_n9509 0.012882f
C6013 a_25860_n9032 a_25559_n10980 0.031194f
C6014 a_26383_1944 VDD 0.559395f
C6015 a_30808_n6334 VDD 0.373881f
C6016 a_26547_n12951 a_26563_n12212 0.08515f
C6017 a_24965_n9860 a_24233_n13388 0.023169f
C6018 a_38380_n11077 a_38292_n10980 0.285629f
C6019 a_43980_n9509 VDD 0.31896f
C6020 a_41292_n12645 a_41740_n12645 0.012882f
C6021 a_37708_n12645 VDD 0.322617f
C6022 a_37484_n15781 VDD 0.322148f
C6023 a_27709_n16132 a_23564_n17700 0.089178f
C6024 a_31324_n4372 a_29744_1564 0.061706f
C6025 a_28300_n18917 VDD 0.329708f
C6026 a_33452_n17349 a_33812_n17252 0.087066f
C6027 a_31436_n18917 a_31884_n18917 0.012882f
C6028 a_45772_n6373 a_46132_n6276 0.087066f
C6029 a_44004_n20008 a_43644_n20052 0.087066f
C6030 a_29532_n10311 a_32543_n9032 0.068784f
C6031 a_28048_1248 VDD 0.022335f
C6032 a_47924_n6276 VDD 0.21239f
C6033 a_41204_n10980 a_41652_n10980 0.013276f
C6034 a_22568_n10512 VDD 0.362677f
C6035 a_43532_n12645 a_43444_n12548 0.285629f
C6036 a_42100_n12548 VDD 0.205948f
C6037 a_32636_n2020 a_33999_n1400 0.013959f
C6038 a_47564_n14213 a_48012_n14213 0.012882f
C6039 a_39276_n14213 a_39188_n14116 0.285629f
C6040 a_42100_n15684 VDD 0.205948f
C6041 a_22052_n4708 a_37585_n3140 0.040578f
C6042 a_43084_n15781 a_43444_n15684 0.087066f
C6043 a_22948_n18820 VDD 0.205626f
C6044 a_30092_1564 a_30296_1564 0.048436f
C6045 a_30604_1515 a_30500_1564 0.026665f
C6046 a_29744_1564 a_31961_1204 0.020455f
C6047 a_33812_n17252 a_34260_n17252 0.013276f
C6048 a_39164_n4805 a_39076_n4708 0.285629f
C6049 a_44428_n17349 a_44340_n17252 0.285629f
C6050 a_29196_n18917 a_29108_n18820 0.285629f
C6051 a_43444_n7844 a_43556_n9032 0.026657f
C6052 a_47452_n20052 a_47900_n20052 0.012001f
C6053 a_27281_n16854 a_24964_n14116 0.023808f
C6054 a_25573_n12167 a_24152_n11680 0.015112f
C6055 a_26861_n10135 a_27485_n10068 0.104193f
C6056 a_39524_n7464 VDD 0.210243f
C6057 a_22352_n12097 a_24464_n11680 0.277491f
C6058 a_22264_n8988 a_22140_n15348 0.080258f
C6059 a_37284_n10600 VDD 0.232632f
C6060 a_45236_n12548 a_45684_n12548 0.013276f
C6061 a_30903_n13780 VDD 1.37524f
C6062 a_27988_n4328 a_22820_n2804 0.042712f
C6063 a_44316_n1669 a_44764_n1669 0.013103f
C6064 a_35716_n16872 VDD 0.207033f
C6065 a_45236_n15684 a_45684_n15684 0.013276f
C6066 a_45324_n3237 a_45684_n3140 0.087066f
C6067 a_44788_n18820 VDD 0.225489f
C6068 a_43892_n4708 a_44340_n4708 0.013276f
C6069 a_32455_n7420 a_32351_n7376 0.277491f
C6070 a_26420_n18820 a_26868_n18820 0.013276f
C6071 a_39724_n18917 a_40084_n18820 0.087066f
C6072 a_24492_n5156 a_28624_n9394 0.068462f
C6073 a_45772_n101 a_46220_n101 0.012552f
C6074 a_39972_n4328 VDD 0.207813f
C6075 a_28435_n10599 a_30808_n10600 0.013167f
C6076 a_32732_n10556 a_32424_n10512 0.934191f
C6077 a_26643_n8292 VDD 0.319115f
C6078 a_36164_n12168 a_36612_n12168 0.013276f
C6079 a_47900_n10644 VDD 0.335152f
C6080 a_40652_n1572 a_45236_n4 0.020613f
C6081 a_40956_n13780 VDD 0.330158f
C6082 a_23608_n15260 a_23912_n15216 0.031502f
C6083 a_22948_n14820 a_25160_n14816 0.042802f
C6084 a_44004_n1192 a_44228_n1192 0.138212f
C6085 a_42748_n16916 VDD 0.315469f
C6086 a_21604_n3844 a_23816_n3840 0.042802f
C6087 a_22364_n4240 a_22568_n4240 0.048436f
C6088 a_22016_n4257 a_24233_n3980 0.020455f
C6089 a_30340_n20008 VDD 0.210296f
C6090 a_24233_n5548 a_24128_n5408 0.116059f
C6091 a_25188_n18440 a_25276_n18484 0.285629f
C6092 a_21692_n18484 a_22140_n18484 0.013103f
C6093 a_39076_n7464 a_39164_n7508 0.285629f
C6094 a_26719_n7464 a_26973_n8292 0.010697f
C6095 a_42660_n7464 a_43108_n7464 0.013276f
C6096 a_44316_n1236 VDD 0.324809f
C6097 a_35804_n20485 a_36164_n20388 0.087174f
C6098 a_46780_n20485 a_47228_n20485 0.013103f
C6099 a_43556_n9032 a_43644_n9076 0.285629f
C6100 a_40420_n10600 a_40868_n10600 0.013276f
C6101 a_47197_908 VDD 0.689874f
C6102 a_42636_n11077 VDD 0.313885f
C6103 a_21604_n708 a_22876_n1148 0.05539f
C6104 a_33452_n14213 VDD 0.301903f
C6105 a_33812_n15304 a_33900_n15348 0.285629f
C6106 a_22672_n2759 a_23319_n2759 0.068833f
C6107 a_25547_n2445 a_25895_n2624 0.317251f
C6108 a_22820_n2804 a_27628_n3841 0.029581f
C6109 a_27988_n4328 a_25237_n4327 1.08764f
C6110 a_40172_n17349 VDD 0.315469f
C6111 a_32220_n16916 a_32668_n16916 0.013103f
C6112 a_35716_n16872 a_35804_n16916 0.285629f
C6113 a_22052_n4708 a_26154_n4536 0.012354f
C6114 a_28492_332 a_32579_769 0.21223f
C6115 a_44004_n20008 VDD 0.2108f
C6116 a_24672_n11339 a_24264_n6976 0.030991f
C6117 a_24492_n5156 a_26095_n7464 0.01417f
C6118 a_23479_n5156 a_26943_n7442 0.25381f
C6119 a_22220_n9860 a_22464_n7393 0.023711f
C6120 a_29892_n18440 a_29532_n18484 0.087066f
C6121 a_47228_n20485 a_47140_n20388 0.285629f
C6122 a_47004_n9076 a_47452_n9076 0.012222f
C6123 a_41740_n4805 VDD 0.313885f
C6124 a_41404_n12212 a_41852_n12212 0.012882f
C6125 a_21940_n11684 VDD 1.84441f
C6126 a_37732_n13736 a_37372_n13780 0.087066f
C6127 a_29444_n708 a_30716_n1148 0.05539f
C6128 a_37844_n14116 VDD 0.214349f
C6129 a_46916_n1572 a_46916_n2760 0.05841f
C6130 a_41316_n15304 a_41764_n15304 0.013276f
C6131 a_32432_n2689 a_34649_n2412 0.020455f
C6132 a_37732_n15304 a_37820_n15348 0.285629f
C6133 a_41204_n17252 VDD 0.226701f
C6134 a_39524_n16872 a_39164_n16916 0.087066f
C6135 a_43108_n4328 a_43556_n4328 0.013276f
C6136 a_39524_n4328 a_39164_n4372 0.087174f
C6137 a_35119_398 a_30104_n1148 0.019491f
C6138 a_31996_n20485 VDD 0.336653f
C6139 a_36252_n18484 a_36700_n18484 0.012001f
C6140 a_27988_n4328 a_28927_n10160 0.031809f
C6141 a_26980_n20008 a_26620_n20052 0.087066f
C6142 a_44092_n7508 a_43980_n7941 0.026339f
C6143 a_25685_n7463 a_25860_n9032 0.012201f
C6144 a_25573_n12167 a_27485_n10068 0.477372f
C6145 a_47140_n20388 a_47588_n20388 0.013276f
C6146 a_22264_n5852 VDD 0.461256f
C6147 a_34652_n11391 a_34538_n10980 0.01244f
C6148 a_23564_n11428 a_24684_n16432 0.039415f
C6149 a_34895_376 a_35156_n325 0.010232f
C6150 a_44004_n9032 VDD 0.2108f
C6151 a_35804_n12212 VDD 0.313975f
C6152 a_44092_n13780 a_44540_n13780 0.012001f
C6153 a_33364_n15304 VDD 0.203482f
C6154 a_27628_n3841 a_25237_n4327 0.151661f
C6155 a_35692_n15348 a_35692_n15781 0.05841f
C6156 a_41988_n2760 a_41628_n2804 0.087174f
C6157 a_31324_n4372 a_31392_n2760 0.014618f
C6158 a_29892_n18440 VDD 0.209775f
C6159 a_46020_n16872 a_46468_n16872 0.013276f
C6160 a_40776_770 a_40260_n408 0.903702f
C6161 a_39544_420 a_40672_864 0.048436f
C6162 a_32356_n20388 VDD 0.214728f
C6163 a_43556_n18440 a_43196_n18484 0.087066f
C6164 a_33476_n20008 a_33924_n20008 0.013276f
C6165 a_29892_n20008 a_29980_n20052 0.285629f
C6166 a_40172_n5940 VDD 0.329275f
C6167 a_30871_n11728 a_32026_n12168 0.037134f
C6168 a_45212_n12212 a_45324_n12645 0.026339f
C6169 a_45660_n12212 VDD 0.320877f
C6170 a_40508_n13780 a_40620_n14213 0.026339f
C6171 a_46468_n1192 a_46556_n1236 0.285629f
C6172 a_40956_n15348 VDD 0.330158f
C6173 a_22052_n15684 a_22500_n15684 0.013276f
C6174 a_42748_n15348 a_42636_n15781 0.026339f
C6175 a_47812_n2760 a_47452_n2804 0.086635f
C6176 a_42604_n2020 a_46556_n1236 0.012909f
C6177 a_31076_376 a_33999_n1400 0.013234f
C6178 a_43556_n18440 VDD 0.209225f
C6179 a_40060_n4372 a_40060_n4805 0.05841f
C6180 a_25530_n5112 a_26154_n4536 0.107109f
C6181 a_23887_n5156 a_22220_n9860 0.03307f
C6182 a_22544_n4690 a_22564_n5112 0.569757f
C6183 a_47004_n18484 a_47452_n18484 0.012222f
C6184 a_35916_n4 VDD 0.010384f
C6185 a_38516_n7844 a_38964_n7844 0.013276f
C6186 a_45772_n7941 a_46132_n7844 0.087066f
C6187 a_45572_n2760 VDD 0.210857f
C6188 a_27302_n9816 a_27485_n10068 0.034561f
C6189 a_25759_1944 VDD 0.723894f
C6190 a_39276_n9509 a_39636_n9412 0.087174f
C6191 a_30215_n6265 VDD 0.824281f
C6192 a_21772_n9860 a_26470_n13736 0.067917f
C6193 a_24684_n16432 a_22600_n12124 0.476633f
C6194 a_24964_n14116 a_26563_n12212 0.020606f
C6195 a_45772_n11077 a_46220_n11077 0.012882f
C6196 a_37932_n11077 a_38292_n10980 0.087174f
C6197 a_43532_n9509 VDD 0.317216f
C6198 a_37260_n12645 VDD 0.31985f
C6199 a_36588_n14213 a_37036_n14213 0.012882f
C6200 a_37036_n15781 VDD 0.334604f
C6201 a_25600_n5895 a_28583_n3140 0.07162f
C6202 a_43868_n2804 a_43980_n3237 0.026339f
C6203 a_28736_1944 a_28836_376 0.417859f
C6204 a_25084_1564 a_29332_1243 0.020443f
C6205 a_47364_1944 a_47452_1900 0.285629f
C6206 a_27852_n18917 VDD 0.329651f
C6207 a_43532_n17349 a_43980_n17349 0.012882f
C6208 a_33452_n17349 a_33364_n17252 0.285629f
C6209 a_22220_n9860 a_22772_n8944 0.024554f
C6210 a_45772_n6373 a_45684_n6276 0.285629f
C6211 a_39860_n6276 a_40308_n6276 0.013276f
C6212 a_39612_n20052 a_40060_n20052 0.012882f
C6213 a_29532_n10311 a_31919_n9032 0.021629f
C6214 a_43556_n20008 a_43644_n20052 0.285629f
C6215 a_36112_n3456 VDD 0.022335f
C6216 a_42548_n9412 a_42996_n9412 0.013276f
C6217 a_28153_1204 VDD 0.480012f
C6218 a_47476_n6276 VDD 0.206217f
C6219 a_34350_n10980 a_35268_n12168 0.012918f
C6220 a_22364_n10512 VDD 0.010384f
C6221 a_34036_n12548 a_34484_n12548 0.013276f
C6222 a_43084_n12645 a_43444_n12548 0.087066f
C6223 a_41652_n12548 VDD 0.205948f
C6224 a_33375_n1976 a_32308_n1976 0.033729f
C6225 a_38828_n14213 a_39188_n14116 0.087066f
C6226 a_41652_n15684 VDD 0.205948f
C6227 a_43084_n15781 a_42996_n15684 0.285629f
C6228 a_34260_n15684 a_34708_n15684 0.013276f
C6229 a_42604_n2020 a_46020_n1572 0.015294f
C6230 a_30604_1515 a_30296_1564 0.934191f
C6231 a_29744_1564 a_31544_1248 0.510371f
C6232 a_22500_n18820 VDD 0.203482f
C6233 a_38716_n4805 a_39076_n4708 0.086905f
C6234 a_43980_n17349 a_44340_n17252 0.087066f
C6235 a_44876_n4805 a_45324_n4805 0.012882f
C6236 a_42188_n18917 a_42636_n18917 0.012882f
C6237 a_28748_n18917 a_29108_n18820 0.087066f
C6238 a_23324_n7420 a_24264_n6976 0.056721f
C6239 a_37820_n20052 a_37820_n20485 0.05841f
C6240 a_47924_n3140 VDD 0.21239f
C6241 a_40652_n1572 VDD 1.77317f
C6242 a_25020_n11383 a_33900_n11428 0.256061f
C6243 a_25573_n12167 a_24569_n11820 0.142814f
C6244 a_23816_n10112 a_24128_n10112 0.119687f
C6245 a_39076_n7464 VDD 0.213966f
C6246 a_47028_n4 a_46916_n1192 0.026657f
C6247 a_36388_n1572 a_34953_n1572 0.036541f
C6248 a_41204_n14116 a_41652_n14116 0.013276f
C6249 a_35268_n16872 VDD 0.207033f
C6250 a_25237_n4327 a_36520_n3868 0.012821f
C6251 a_45324_n3237 a_45236_n3140 0.285629f
C6252 a_44340_n18820 VDD 0.212826f
C6253 a_44340_n17252 a_44788_n17252 0.013276f
C6254 a_39724_n18917 a_39636_n18820 0.285629f
C6255 a_29123_n6679 a_31965_n8292 0.472234f
C6256 a_32455_n7420 a_33048_n7420 0.361958f
C6257 a_31799_n7508 a_32856_n7376 0.056721f
C6258 a_22772_n1104 VDD 0.298894f
C6259 a_35356_n20485 a_35804_n20485 0.013103f
C6260 a_39524_n4328 VDD 0.210243f
C6261 a_31872_n10529 a_32424_n10512 0.361958f
C6262 a_24752_n8292 VDD 0.584827f
C6263 a_29540_n11728 a_30180_n12168 0.010102f
C6264 a_31279_n11728 a_30599_n12167 0.190494f
C6265 a_47452_n10644 VDD 0.313885f
C6266 a_37620_n12548 a_37732_n13736 0.026657f
C6267 a_43644_n705 a_47564_n101 0.029694f
C6268 a_42772_n4 a_42884_n1192 0.026657f
C6269 a_40508_n13780 VDD 0.313885f
C6270 a_23360_n15233 a_23912_n15216 0.361958f
C6271 a_22948_n14820 a_25577_n14956 0.019043f
C6272 a_23608_n15260 a_23708_n15216 0.092638f
C6273 a_44228_n1572 a_44676_n1572 0.013276f
C6274 a_42300_n16916 VDD 0.315469f
C6275 a_22876_n4284 a_22568_n4240 0.934191f
C6276 a_38740_n15684 a_38628_n16872 0.026657f
C6277 a_21604_n3844 a_24233_n3980 0.019043f
C6278 a_29892_n20008 VDD 0.208807f
C6279 a_44004_n1192 a_40260_n408 0.084018f
C6280 a_25188_n18440 a_24828_n18484 0.086742f
C6281 a_22948_n18820 a_22948_n20008 0.05841f
C6282 a_39076_n7464 a_38716_n7508 0.087066f
C6283 a_36948_n18820 a_37396_n18820 0.013276f
C6284 a_35804_n20485 a_35716_n20388 0.285629f
C6285 a_39164_n9076 a_39612_n9076 0.012882f
C6286 a_43556_n9032 a_43196_n9076 0.087066f
C6287 a_29532_n10311 a_28335_n10644 0.856216f
C6288 a_25573_n12167 a_27526_n9816 0.066157f
C6289 a_22544_n4690 VDD 0.537892f
C6290 a_23564_n8292 a_22016_n13665 0.027741f
C6291 a_26861_n10135 a_26543_n11384 0.03239f
C6292 a_46573_841 VDD 0.571865f
C6293 a_39076_n12168 a_39524_n12168 0.013276f
C6294 a_42188_n11077 VDD 0.313885f
C6295 a_32413_n14564 VDD 0.769827f
C6296 a_24771_n2804 a_25895_n2624 0.152869f
C6297 a_33812_n15304 a_33452_n15348 0.087174f
C6298 a_25547_n2445 a_26499_n2732 0.869605f
C6299 a_39724_n17349 VDD 0.318714f
C6300 a_35716_n16872 a_35356_n16916 0.086742f
C6301 a_22052_n4708 a_25530_n5112 0.014671f
C6302 a_45684_n15684 a_45572_n16872 0.026657f
C6303 a_43556_n20008 VDD 0.209225f
C6304 a_29444_n18440 a_29532_n18484 0.285629f
C6305 a_39357_n5364 a_40084_n5896 0.169527f
C6306 a_23479_n5156 a_26719_n7464 0.046723f
C6307 a_33028_n18440 a_33476_n18440 0.013276f
C6308 a_24492_n5156 a_25685_n7463 0.035784f
C6309 a_22220_n9860 a_22052_n6980 0.013023f
C6310 a_24672_n11339 a_24681_n7116 0.041412f
C6311 a_27988_n4328 a_25020_n11383 0.352323f
C6312 a_45572_n7464 a_46020_n7464 0.013276f
C6313 a_30004_n18820 a_29892_n20008 0.026657f
C6314 a_25972_n6276 a_28225_n9031 0.090796f
C6315 a_23479_n5156 a_26239_n11428 0.048464f
C6316 VDD XRST 0.265981f
C6317 a_31348_n1931 VDD 0.455129f
C6318 a_46780_n20485 a_47140_n20388 0.087174f
C6319 a_35716_n20388 a_36164_n20388 0.013276f
C6320 a_41292_n4805 VDD 0.31945f
C6321 a_43196_n10644 a_43644_n10644 0.012882f
C6322 a_21872_n9394 VDD 0.538427f
C6323 a_32026_n12168 a_32413_n12996 0.033256f
C6324 a_34068_n4 a_34271_n1192 0.043031f
C6325 a_47924_n10980 VDD 0.21239f
C6326 a_40868_n13736 a_41316_n13736 0.013276f
C6327 a_29444_n708 a_29856_n1121 0.536965f
C6328 a_37284_n13736 a_37372_n13780 0.285629f
C6329 a_37396_n14116 VDD 0.211702f
C6330 a_32780_n2672 a_32984_n2672 0.048436f
C6331 a_37732_n15304 a_37372_n15348 0.087066f
C6332 a_40532_n17252 VDD 0.212412f
C6333 a_39076_n4328 a_39164_n4372 0.285629f
C6334 a_39076_n16872 a_39164_n16916 0.285629f
C6335 a_42660_n16872 a_43108_n16872 0.013276f
C6336 a_34895_376 a_30104_n1148 0.024826f
C6337 a_31548_n20485 VDD 0.360143f
C6338 a_43308_n5940 a_43756_n5940 0.012222f
C6339 a_27988_n4328 a_28437_n13705 0.034789f
C6340 a_22588_n20052 a_23036_n20052 0.012882f
C6341 a_26532_n20008 a_26620_n20052 0.285629f
C6342 a_27302_n9816 a_27526_n9816 0.75472f
C6343 a_25573_n12167 a_26861_n10135 0.081307f
C6344 a_43196_n9076 a_43084_n9509 0.026339f
C6345 a_25237_n10599 a_22220_n12996 0.045365f
C6346 a_22016_n5825 VDD 0.800064f
C6347 a_39164_n10644 a_39276_n11077 0.026339f
C6348 a_43556_n9032 VDD 0.209225f
C6349 a_35356_n12212 VDD 0.317587f
C6350 a_23816_n704 a_24578_n2020 0.023779f
C6351 a_41203_n799 a_41533_n727 0.538085f
C6352 a_32916_n15304 VDD 0.172738f
C6353 a_44092_n15348 a_44540_n15348 0.012001f
C6354 a_41540_n2760 a_41628_n2804 0.285629f
C6355 a_31324_n4372 a_31412_n2276 0.040431f
C6356 a_29444_n18440 VDD 0.229103f
C6357 a_45572_n4328 a_46020_n4328 0.013276f
C6358 a_42771_769 a_43101_841 0.538085f
C6359 a_38951_420 a_40672_864 0.401636f
C6360 a_31908_n20388 VDD 0.211263f
C6361 a_39164_n18484 a_39612_n18484 0.012882f
C6362 a_43108_n18440 a_43196_n18484 0.285629f
C6363 a_29892_n20008 a_29532_n20052 0.087066f
C6364 a_41740_n7941 a_42188_n7941 0.012882f
C6365 a_30871_n11728 a_31279_n11728 0.044274f
C6366 a_28232_n12606 a_29360_n12864 0.048436f
C6367 a_45212_n12212 VDD 0.342281f
C6368 a_26532_n14437 a_27496_n14116 0.08126f
C6369 a_46468_n1192 a_46108_n1236 0.086905f
C6370 a_40508_n15348 VDD 0.313885f
C6371 a_45660_n2804 a_46108_n2804 0.012552f
C6372 a_47364_n2760 a_47452_n2804 0.285629f
C6373 a_42604_n2020 a_46108_n1236 0.052966f
C6374 a_43108_n18440 VDD 0.206217f
C6375 a_32108_n17349 a_32556_n17349 0.012001f
C6376 a_23479_n5156 a_22220_n9860 0.277319f
C6377 a_25237_n5895 a_26154_n4536 0.054242f
C6378 a_39500_n6373 a_39948_n6373 0.012222f
C6379 a_41204_1243 OUT[4] 0.016632f
C6380 a_36428_n53 VDD 0.248737f
C6381 a_36252_n20052 a_36700_n20052 0.012001f
C6382 a_45772_n7941 a_45684_n7844 0.285629f
C6383 a_45124_n2760 VDD 0.260375f
C6384 a_39276_n9509 a_39188_n9412 0.285629f
C6385 a_46668_n9509 a_47116_n9509 0.012882f
C6386 a_37932_n11077 a_37844_n10980 0.285629f
C6387 a_21772_n9860 a_26266_n13736 0.038529f
C6388 a_43084_n9509 VDD 0.313885f
C6389 a_36812_n12645 VDD 0.319488f
C6390 a_36588_n15781 VDD 0.299665f
C6391 a_40172_n15781 a_40620_n15781 0.012001f
C6392 a_23564_n20836 a_23564_n17700 0.106598f
C6393 a_22164_n2760 a_28225_n4327 0.087046f
C6394 a_23004_n2332 a_22672_n2759 0.108617f
C6395 a_24631_n3588 a_23507_n2759 0.038903f
C6396 a_27404_n18917 VDD 0.329651f
C6397 a_24492_n5156 a_28617_n8548 0.44043f
C6398 a_30988_n18917 a_31436_n18917 0.012882f
C6399 a_45324_n6373 a_45684_n6276 0.087066f
C6400 a_43556_n20008 a_43196_n20052 0.087066f
C6401 a_23479_n5156 a_27279_n12146 0.067347f
C6402 a_36217_n3500 VDD 0.483571f
C6403 a_32581_n9860 a_32424_n10512 0.056633f
C6404 a_27736_1248 VDD 1.33472f
C6405 a_47028_n6276 VDD 0.206217f
C6406 a_22876_n10556 VDD 0.248203f
C6407 a_43084_n12645 a_42996_n12548 0.285629f
C6408 a_41204_n12548 VDD 0.227793f
C6409 a_32860_n2020 a_32308_n1976 0.014392f
C6410 a_47116_n14213 a_47564_n14213 0.012882f
C6411 a_38828_n14213 a_38740_n14116 0.285629f
C6412 a_41204_n15684 VDD 0.226701f
C6413 a_23564_n20836 a_23932_n16916 0.04507f
C6414 a_42636_n15781 a_42996_n15684 0.087066f
C6415 a_22052_n18820 VDD 0.203482f
C6416 a_38716_n4805 a_38628_n4708 0.285629f
C6417 a_43980_n17349 a_43892_n17252 0.285629f
C6418 a_33364_n17252 a_33812_n17252 0.013276f
C6419 a_23228_n6679 a_22568_n5808 0.019564f
C6420 a_28748_n18917 a_28660_n18820 0.285629f
C6421 a_42996_n7844 a_43108_n9032 0.026657f
C6422 a_47004_n20052 a_47452_n20052 0.012222f
C6423 a_47476_n3140 VDD 0.206217f
C6424 a_26531_n10207 a_26861_n10135 0.538085f
C6425 a_24233_n10252 a_24128_n10112 0.116059f
C6426 a_25860_n9032 a_26563_n12212 0.013524f
C6427 a_25020_n11383 a_34652_n11391 0.108469f
C6428 a_45100_1467 VDD 0.354119f
C6429 a_38628_n7464 VDD 0.214f
C6430 a_23564_n11428 a_23949_n12996 0.019613f
C6431 a_21772_n9860 a_26532_n14437 0.048714f
C6432 a_24964_n14116 a_21872_n12530 0.033725f
C6433 a_33900_n11428 VDD 0.722913f
C6434 a_44788_n12548 a_45236_n12548 0.013276f
C6435 a_35816_n174 a_35916_n4 0.083421f
C6436 a_27820_n16432 VDD 0.649674f
C6437 a_43868_n1669 a_44316_n1669 0.013103f
C6438 a_34820_n16872 VDD 0.207033f
C6439 a_44876_n3237 a_45236_n3140 0.087066f
C6440 a_44788_n15684 a_45236_n15684 0.013276f
C6441 a_25237_n4327 a_35848_n3868 0.494265f
C6442 a_43892_n18820 VDD 0.210221f
C6443 a_43444_n4708 a_43892_n4708 0.013276f
C6444 a_32560_n7020 a_33048_n7420 0.08126f
C6445 a_29123_n6679 a_31341_n8292 0.067685f
C6446 a_39276_n18917 a_39636_n18820 0.087066f
C6447 a_24492_n5156 a_27281_n16854 0.649154f
C6448 a_22220_n9860 a_21892_n9816 0.526558f
C6449 a_25972_n18820 a_26420_n18820 0.013276f
C6450 a_24128_n704 VDD 0.022903f
C6451 a_45324_n101 a_45772_n101 0.012552f
C6452 a_39076_n4328 VDD 0.14097f
C6453 a_31460_n10116 a_33672_n10112 0.042802f
C6454 a_31872_n10529 a_32220_n10512 0.401636f
C6455 a_23564_n8292 VDD 1.4269f
C6456 a_35716_n12168 a_36164_n12168 0.013276f
C6457 a_32026_n12168 a_31760_n12168 0.128352f
C6458 a_47004_n10644 VDD 0.313885f
C6459 a_40060_n13780 VDD 0.314419f
C6460 a_23360_n15233 a_23708_n15216 0.401636f
C6461 a_27192_n14286 a_26755_n16132 0.050006f
C6462 a_23608_n15260 a_24220_n15260 0.042372f
C6463 a_41852_n16916 VDD 0.315469f
C6464 a_44004_n1192 a_43725_908 0.067844f
C6465 a_37859_377 a_39804_464 0.028439f
C6466 a_29444_n20008 VDD 0.226701f
C6467 a_24740_n18440 a_24828_n18484 0.285629f
C6468 a_22568_n5808 a_22772_n5808 0.66083f
C6469 a_38628_n7464 a_38716_n7508 0.285629f
C6470 a_42212_n7464 a_42660_n7464 0.013276f
C6471 a_43556_n661 VDD 0.479342f
C6472 a_25573_n12167 a_27302_n9816 0.058036f
C6473 a_46332_n20485 a_46780_n20485 0.013103f
C6474 a_35356_n20485 a_35716_n20388 0.087174f
C6475 a_43108_n9032 a_43196_n9076 0.285629f
C6476 a_39972_n10600 a_40420_n10600 0.013276f
C6477 a_46243_769 VDD 0.311024f
C6478 a_25573_n12167 a_21772_n12996 0.01998f
C6479 a_41740_n11077 VDD 0.313885f
C6480 a_31789_n14564 VDD 0.576678f
C6481 a_22820_n2804 a_31292_n2804 0.028825f
C6482 a_33364_n15304 a_33452_n15348 0.285629f
C6483 a_23404_816 a_25732_n1192 0.01472f
C6484 a_23004_n2332 a_22016_n1121 0.038594f
C6485 a_39276_n17349 VDD 0.320362f
C6486 a_22052_n4708 a_25237_n5895 0.023286f
C6487 a_31772_n16916 a_32220_n16916 0.013103f
C6488 a_35268_n16872 a_35356_n16916 0.285629f
C6489 a_47924_n4 a_47812_n1192 0.026657f
C6490 a_28492_332 a_24631_n3588 0.037887f
C6491 a_43108_n20008 VDD 0.206217f
C6492 a_47476_n18820 a_47924_n18820 0.013276f
C6493 a_27988_n4328 VDD 1.00058f
C6494 a_46780_n20485 a_46692_n20388 0.285629f
C6495 a_46556_n9076 a_47004_n9076 0.012222f
C6496 a_40508_n4805 VDD 0.318168f
C6497 a_27485_n8500 VDD 0.70259f
C6498 a_24964_n14116 a_29479_n13735 0.076055f
C6499 a_40956_n12212 a_41404_n12212 0.012882f
C6500 a_42604_n2020 a_46668_n101 0.010099f
C6501 a_47476_n10980 VDD 0.206217f
C6502 a_25132_n16432 a_25160_n14816 0.061841f
C6503 a_36948_n14116 VDD 0.21223f
C6504 a_40868_n15304 a_41316_n15304 0.013276f
C6505 a_37284_n15304 a_37372_n15348 0.285629f
C6506 a_33292_n2716 a_32984_n2672 0.934191f
C6507 a_46468_n1572 a_46468_n2760 0.05841f
C6508 a_40084_n17252 VDD 0.206509f
C6509 a_42660_n4328 a_43108_n4328 0.013276f
C6510 a_39076_n16872 a_38716_n16916 0.087066f
C6511 a_31100_n20485 VDD 0.339976f
C6512 a_34271_376 a_30104_n1148 0.021996f
C6513 a_35804_n18484 a_36252_n18484 0.012882f
C6514 a_26532_n20008 a_26172_n20052 0.087066f
C6515 a_43644_n7508 a_43532_n7941 0.026339f
C6516 a_46692_n20388 a_47140_n20388 0.013276f
C6517 a_24965_n9860 a_22220_n12996 0.130062f
C6518 a_25573_n12167 a_26531_n10207 0.030716f
C6519 a_21604_n5412 VDD 1.86146f
C6520 a_26547_n12951 a_26543_n11384 0.469862f
C6521 a_34403_332 a_35156_n325 0.030696f
C6522 a_43108_n9032 VDD 0.206217f
C6523 a_28300_n15348 a_30555_n13780 0.028784f
C6524 a_43644_n13780 a_44092_n13780 0.012882f
C6525 a_35244_n15348 a_35244_n15781 0.05841f
C6526 a_41540_n2760 a_41180_n2804 0.087174f
C6527 a_31324_n4372 a_30555_n2729 0.263546f
C6528 a_28524_n18484 VDD 0.349067f
C6529 a_45572_n16872 a_46020_n16872 0.013276f
C6530 a_31460_n20388 VDD 0.244018f
C6531 a_39056_820 a_40672_864 0.011851f
C6532 a_40776_770 a_43101_841 0.016309f
C6533 a_43108_n18440 a_42748_n18484 0.087066f
C6534 a_29444_n20008 a_29532_n20052 0.285629f
C6535 a_33028_n20008 a_33476_n20008 0.013276f
C6536 a_27628_n3841 VDD 0.548782f
C6537 a_26470_n9322 VDD 0.760321f
C6538 a_27639_n12537 a_29360_n12864 0.401636f
C6539 a_47812_n12168 VDD 0.211703f
C6540 a_40060_n13780 a_40172_n14213 0.026339f
C6541 a_46020_n1192 a_46108_n1236 0.285629f
C6542 a_26532_n14437 a_27292_n14116 0.011851f
C6543 a_47364_n1192 a_47812_n1192 0.013276f
C6544 a_40060_n15348 VDD 0.314419f
C6545 a_21604_n15684 a_22052_n15684 0.013276f
C6546 a_24088_n16087 a_23564_n20836 0.194319f
C6547 a_42300_n15348 a_42188_n15781 0.026339f
C6548 a_47364_n2760 a_47004_n2804 0.086742f
C6549 a_42604_n2020 a_45660_n1236 0.02233f
C6550 a_42660_n18440 VDD 0.206217f
C6551 a_44540_n16916 a_44428_n17349 0.026339f
C6552 a_22444_n5156 a_22564_n5112 0.393749f
C6553 a_39612_n4372 a_39612_n4805 0.05841f
C6554 a_25237_n5895 a_25530_n5112 0.517287f
C6555 a_27988_n4328 a_27167_n10808 0.010341f
C6556 a_46556_n18484 a_47004_n18484 0.012222f
C6557 a_38068_n7844 a_38516_n7844 0.013276f
C6558 a_45324_n7941 a_45684_n7844 0.087066f
C6559 a_44316_n2804 VDD 0.3424f
C6560 a_38828_n9509 a_39188_n9412 0.087174f
C6561 a_22052_1944 VDD 1.2611f
C6562 a_29123_n6679 VDD 1.10117f
C6563 a_37484_n11077 a_37844_n10980 0.087174f
C6564 a_45324_n11077 a_45772_n11077 0.012882f
C6565 a_42636_n9509 VDD 0.313885f
C6566 a_36364_n12645 VDD 0.316395f
C6567 a_36140_n14213 a_36588_n14213 0.012882f
C6568 a_36140_n15781 VDD 0.296789f
C6569 a_43420_n2804 a_43532_n3237 0.026339f
C6570 a_31324_n4372 a_29332_1243 0.015662f
C6571 a_26956_n18917 VDD 0.328067f
C6572 a_43084_n17349 a_43532_n17349 0.012882f
C6573 a_32556_n17349 a_32468_n17252 0.285629f
C6574 a_45324_n6373 a_45236_n6276 0.285629f
C6575 a_25612_n6679 a_31451_n7508 0.013249f
C6576 a_39164_n20052 a_39612_n20052 0.012882f
C6577 a_43108_n20008 a_43196_n20052 0.285629f
C6578 a_23479_n5156 a_27055_n12168 0.056416f
C6579 a_35800_n3456 VDD 1.32948f
C6580 a_42100_n9412 a_42548_n9412 0.013276f
C6581 a_26692_1564 VDD 0.298894f
C6582 a_46580_n6276 VDD 0.209016f
C6583 a_22016_n10529 VDD 0.808133f
C6584 a_28121_n10980 a_27852_n14990 0.362159f
C6585 a_42636_n12645 a_42996_n12548 0.087066f
C6586 a_40308_n12548 VDD 0.212323f
C6587 a_32636_n2020 a_32308_n1976 1.29386f
C6588 a_38380_n14213 a_38740_n14116 0.087066f
C6589 a_40532_n15684 VDD 0.212412f
C6590 a_33812_n15684 a_34260_n15684 0.013276f
C6591 a_42636_n15781 a_42548_n15684 0.285629f
C6592 a_23564_n20836 a_23484_n16916 0.013064f
C6593 a_21604_n18820 VDD 0.221763f
C6594 a_29332_1243 a_31961_1204 0.019043f
C6595 a_28836_376 a_30092_1564 0.088321f
C6596 a_29744_1564 a_30296_1564 0.361958f
C6597 a_44428_n4805 a_44876_n4805 0.012882f
C6598 a_25237_n5895 a_23816_n5408 0.014425f
C6599 a_24492_n5156 a_24128_n5408 0.011361f
C6600 a_38268_n4805 a_38628_n4708 0.086905f
C6601 a_43532_n17349 a_43892_n17252 0.087066f
C6602 a_41740_n18917 a_42188_n18917 0.012882f
C6603 a_28300_n18917 a_28660_n18820 0.087066f
C6604 a_22464_n7393 a_24264_n6976 0.510371f
C6605 a_37372_n20052 a_37372_n20485 0.05841f
C6606 a_47028_n3140 VDD 0.206217f
C6607 a_43728_1248 VDD 0.024223f
C6608 a_38180_n7464 VDD 0.239345f
C6609 a_34652_n11391 VDD 0.981395f
C6610 a_35940_n1931 a_34953_n1572 0.022441f
C6611 a_35288_n1975 a_34248_n3310 0.19494f
C6612 a_34372_n16872 VDD 0.207033f
C6613 a_39860_n3140 a_40308_n3140 0.013276f
C6614 a_44876_n3237 a_44788_n3140 0.285629f
C6615 a_22052_n4708 a_21792_n7464 0.126026f
C6616 a_24631_n3588 a_27932_n3543 0.080079f
C6617 a_43444_n18820 VDD 0.208815f
C6618 a_31324_n4372 a_31076_376 0.027819f
C6619 a_43892_n17252 a_44340_n17252 0.013276f
C6620 a_29123_n6679 a_30676_n7844 0.7031f
C6621 a_32560_n7020 a_32455_n7420 0.536965f
C6622 a_31799_n7508 a_32351_n7376 0.119687f
C6623 a_34068_n4 VDD 0.598557f
C6624 a_39276_n18917 a_39188_n18820 0.285629f
C6625 a_34908_n20485 a_35356_n20485 0.013103f
C6626 a_36520_n3868 VDD 0.538731f
C6627 a_31460_n10116 a_34089_n10252 0.019043f
C6628 a_31872_n10529 a_32732_n10556 0.882105f
C6629 a_35119_398 VDD 0.310107f
C6630 a_29540_n11728 a_30599_n12167 0.026863f
C6631 a_31279_n11728 a_31760_n12168 0.064827f
C6632 a_46556_n10644 VDD 0.31705f
C6633 a_37172_n12548 a_37284_n13736 0.026657f
C6634 a_39612_n13780 VDD 0.317476f
C6635 a_43780_n1572 a_44228_n1572 0.013276f
C6636 a_23360_n15233 a_24220_n15260 0.882105f
C6637 a_41404_n16916 VDD 0.315469f
C6638 a_22016_n4257 a_22568_n4240 0.361958f
C6639 a_21792_n7464 a_22364_n4240 0.088321f
C6640 a_38292_n15684 a_38180_n16872 0.026657f
C6641 a_44004_n1192 a_43101_841 0.012916f
C6642 a_28860_n20052 VDD 0.356617f
C6643 a_24740_n18440 a_24380_n18484 0.087174f
C6644 a_24233_n5548 a_23816_n5408 0.633318f
C6645 a_36500_n18820 a_36948_n18820 0.013276f
C6646 a_22500_n18820 a_22500_n20008 0.05841f
C6647 a_26095_n7464 a_26643_n8292 0.017184f
C6648 a_38628_n7464 a_38268_n7508 0.087066f
C6649 a_42972_n1236 VDD 0.321474f
C6650 a_43108_n9032 a_42748_n9076 0.087066f
C6651 a_38716_n9076 a_39164_n9076 0.012882f
C6652 a_34092_n9076 a_34986_n9032 0.02845f
C6653 a_35356_n20485 a_35268_n20388 0.285629f
C6654 a_22444_n5156 VDD 1.42314f
C6655 a_45572_376 VDD 0.208834f
C6656 a_48012_n7941 VDD 0.343411f
C6657 a_22600_n12124 a_22264_n13692 0.11996f
C6658 a_38628_n12168 a_39076_n12168 0.013276f
C6659 a_28300_n15348 a_34572_n12645 0.049052f
C6660 a_41292_n11077 VDD 0.318502f
C6661 a_21604_n708 a_22016_n1121 0.536965f
C6662 a_28752_n15348 VDD 1.21949f
C6663 a_36052_n15304 a_36500_n15304 0.013276f
C6664 a_33364_n15304 a_33004_n15348 0.087174f
C6665 a_38828_n17349 VDD 0.322604f
C6666 a_45236_n15684 a_45124_n16872 0.026657f
C6667 a_35268_n16872 a_34908_n16916 0.086905f
C6668 a_22052_n4708 a_24672_n11339 0.019815f
C6669 a_28492_332 a_30372_376 0.017171f
C6670 a_42660_n20008 VDD 0.206217f
C6671 a_36773_n5468 a_37820_n5940 0.075345f
C6672 a_23479_n5156 a_25685_n7463 0.077623f
C6673 a_32580_n18440 a_33028_n18440 0.013276f
C6674 a_29556_n18820 a_29444_n20008 0.026657f
C6675 a_25612_n6679 a_34092_n9076 0.031511f
C6676 a_45124_n7464 a_45572_n7464 0.013276f
C6677 a_35268_n20388 a_35716_n20388 0.013276f
C6678 a_46332_n20485 a_46692_n20388 0.087174f
C6679 a_40060_n4805 VDD 0.297323f
C6680 a_42748_n10644 a_43196_n10644 0.012882f
C6681 a_26861_n8567 VDD 0.576471f
C6682 a_31279_n11728 a_31789_n12996 0.014021f
C6683 a_47028_n10980 VDD 0.206217f
C6684 a_42604_n2020 a_46220_n101 0.04138f
C6685 a_40420_n13736 a_40868_n13736 0.013276f
C6686 a_36500_n14116 VDD 0.205016f
C6687 a_32432_n2689 a_32984_n2672 0.361958f
C6688 a_24631_n3588 a_30612_n1104 0.011021f
C6689 a_39636_n17252 VDD 0.209407f
C6690 a_38628_n16872 a_38716_n16916 0.285629f
C6691 a_42212_n16872 a_42660_n16872 0.013276f
C6692 a_34403_332 a_30104_n1148 0.034369f
C6693 a_30652_n20485 VDD 0.335905f
C6694 a_42860_n5940 a_43308_n5940 0.013103f
C6695 a_22140_n20052 a_22588_n20052 0.012882f
C6696 a_26084_n20008 a_26172_n20052 0.285629f
C6697 a_34248_n3310 VDD 0.364719f
C6698 a_42748_n9076 a_42636_n9509 0.026339f
C6699 a_21772_n9860 a_25724_n14564 0.024109f
C6700 a_24573_n9860 a_22220_n12996 0.012026f
C6701 a_25573_n12167 a_25412_n10600 0.025285f
C6702 a_38716_n10644 a_38828_n11077 0.026339f
C6703 a_42660_n9032 VDD 0.206217f
C6704 a_28300_n15348 a_30159_n13296 0.024576f
C6705 a_27316_n14820 VDD 0.81684f
C6706 a_43644_n15348 a_44092_n15348 0.012882f
C6707 a_41092_n2760 a_41180_n2804 0.285629f
C6708 a_28076_n18484 VDD 0.329378f
C6709 a_45124_n4328 a_45572_n4328 0.013276f
C6710 a_40260_n408 a_39556_n4 0.223801f
C6711 a_31012_n20388 VDD 0.211403f
C6712 a_40776_770 a_42771_769 0.212887f
C6713 a_44004_n1192 OUT[4] 0.012528f
C6714 a_42660_n18440 a_42748_n18484 0.285629f
C6715 a_38716_n18484 a_39164_n18484 0.012882f
C6716 a_41292_n7941 a_41740_n7941 0.012882f
C6717 a_32020_n2276 VDD 1.80079f
C6718 a_47900_n10644 a_48012_n11077 0.026339f
C6719 a_26266_n9240 VDD 0.597903f
C6720 a_28121_n10980 a_29161_n14476 0.050728f
C6721 a_47364_n12168 VDD 0.205948f
C6722 a_46020_n1192 a_45660_n1236 0.086905f
C6723 a_26532_n14437 a_27804_n14165 0.05539f
C6724 a_39612_n15348 VDD 0.317476f
C6725 a_45212_n2804 a_45660_n2804 0.012552f
C6726 a_46916_n2760 a_47004_n2804 0.285629f
C6727 a_42212_n18440 VDD 0.206217f
C6728 a_22544_n4690 a_22220_n9860 0.064129f
C6729 a_23479_n5156 a_23228_n6679 0.530856f
C6730 a_23887_n5156 a_23207_n4708 0.152057f
C6731 a_31660_n17349 a_32108_n17349 0.012222f
C6732 a_45324_n7941 a_45236_n7844 0.285629f
C6733 a_35804_n20052 a_36252_n20052 0.012882f
C6734 a_43868_n2804 VDD 0.318926f
C6735 a_21604_2475 VDD 0.54595f
C6736 a_25573_n12167 a_24964_n14116 0.969746f
C6737 a_46220_n9509 a_46668_n9509 0.012882f
C6738 a_38828_n9509 a_38740_n9412 0.285629f
C6739 a_30320_n6636 VDD 1.77236f
C6740 a_37484_n11077 a_37396_n10980 0.285629f
C6741 a_42188_n9509 VDD 0.313885f
C6742 a_39948_n12645 a_40396_n12645 0.012001f
C6743 a_35916_n12645 VDD 0.315889f
C6744 a_42157_n660 a_41684_n1976 0.030473f
C6745 a_35692_n15781 VDD 0.296789f
C6746 a_39724_n15781 a_40172_n15781 0.012882f
C6747 a_25084_1564 a_27736_1248 0.027465f
C6748 a_26508_n18917 VDD 0.328067f
C6749 a_32108_n17349 a_32468_n17252 0.086635f
C6750 a_22220_n9860 a_21872_n9394 0.52715f
C6751 a_44876_n6373 a_45236_n6276 0.087066f
C6752 a_30540_n18917 a_30988_n18917 0.012882f
C6753 a_23479_n5156 a_26431_n12168 0.018445f
C6754 a_43108_n20008 a_42748_n20052 0.087066f
C6755 a_34756_n3140 VDD 0.298894f
C6756 a_26488_1564 VDD 0.360598f
C6757 a_32581_n9860 a_32732_n10556 0.015944f
C6758 a_46132_n6276 VDD 0.210512f
C6759 a_40084_n10980 a_40532_n10980 0.013276f
C6760 a_21604_n10116 VDD 1.79673f
C6761 a_42636_n12645 a_42548_n12548 0.285629f
C6762 a_39860_n12548 VDD 0.209112f
C6763 a_38380_n14213 a_38292_n14116 0.285629f
C6764 a_46668_n14213 a_47116_n14213 0.012882f
C6765 a_40084_n15684 VDD 0.206509f
C6766 a_42188_n15781 a_42548_n15684 0.087066f
C6767 a_29332_1243 a_31544_1248 0.042802f
C6768 a_29744_1564 a_30092_1564 0.401636f
C6769 a_48012_n18917 VDD 0.343411f
C6770 a_23228_n6679 a_22876_n5852 0.023921f
C6771 a_43532_n17349 a_43444_n17252 0.285629f
C6772 a_25237_n5895 a_24233_n5548 0.113153f
C6773 a_38268_n4805 a_38180_n4708 0.285629f
C6774 a_22464_n7393 a_24681_n7116 0.020455f
C6775 a_22812_n7376 a_23016_n7376 0.048436f
C6776 a_22052_n6980 a_24264_n6976 0.042802f
C6777 a_28300_n18917 a_28212_n18820 0.285629f
C6778 a_46556_n20052 a_47004_n20052 0.012222f
C6779 a_42548_n7844 a_42660_n9032 0.026657f
C6780 a_46580_n3140 VDD 0.209016f
C6781 a_28335_n10644 a_33900_n11428 0.042863f
C6782 a_22568_n10512 a_22772_n10512 0.66083f
C6783 a_43833_1204 VDD 0.478082f
C6784 a_37732_n7464 VDD 0.209811f
C6785 a_23212_n12124 a_24152_n11680 0.056721f
C6786 a_36324_n4 VDD 0.299594f
C6787 a_32628_n10512 VDD 0.300528f
C6788 a_44340_n12548 a_44788_n12548 0.013276f
C6789 a_35288_n1975 a_34953_n1572 0.019958f
C6790 a_43420_n1669 a_43868_n1669 0.013103f
C6791 a_33924_n16872 VDD 0.207033f
C6792 a_44340_n15684 a_44788_n15684 0.013276f
C6793 a_25237_n4327 a_28225_n4327 0.019081f
C6794 a_44428_n3237 a_44788_n3140 0.087066f
C6795 a_22052_n4708 a_22016_n4257 0.012773f
C6796 a_42996_n18820 VDD 0.206098f
C6797 a_42996_n4708 a_43444_n4708 0.013276f
C6798 a_31451_n7508 a_32351_n7376 0.116059f
C6799 a_29123_n6679 a_28972_n8247 0.10592f
C6800 a_23479_n5156 a_27281_n16854 0.12771f
C6801 a_25524_n18820 a_25972_n18820 0.013276f
C6802 a_33508_n408 VDD 0.566777f
C6803 a_30036_n7464 a_30240_n7464 0.033243f
C6804 a_38828_n18917 a_39188_n18820 0.087066f
C6805 a_27279_n1170 VDD 0.322699f
C6806 a_29532_n10311 a_27281_n16854 0.241964f
C6807 a_35848_n3868 VDD 0.44676f
C6808 a_30808_n10116 a_32220_n10512 0.086679f
C6809 a_34895_376 VDD 0.573255f
C6810 a_33308_n7376 VDD 0.298903f
C6811 a_28927_n10160 a_30555_n13780 0.112506f
C6812 a_35268_n12168 a_35716_n12168 0.013276f
C6813 a_46108_n10644 VDD 0.318654f
C6814 a_39164_n13780 VDD 0.319301f
C6815 a_23360_n15233 a_23608_n15260 0.373398f
C6816 a_22948_n14820 a_23912_n15216 0.08126f
C6817 a_40956_n16916 VDD 0.330158f
C6818 a_21604_n3844 a_22568_n4240 0.08126f
C6819 a_22016_n4257 a_22364_n4240 0.401636f
C6820 a_28412_n20052 VDD 0.315469f
C6821 a_27988_n18440 a_28436_n18440 0.013276f
C6822 a_24292_n18440 a_24380_n18484 0.285629f
C6823 a_22876_n5852 a_22772_n5808 0.026665f
C6824 a_42100_n6276 CLK 0.018145f
C6825 a_38180_n7464 a_38268_n7508 0.285629f
C6826 a_41764_n7464 a_42212_n7464 0.013276f
C6827 a_34908_n20485 a_35268_n20388 0.087174f
C6828 a_45884_n20485 a_46332_n20485 0.013103f
C6829 a_42660_n9032 a_42748_n9076 0.285629f
C6830 a_21604_n5067 VDD 0.536321f
C6831 a_39524_n10600 a_39972_n10600 0.013276f
C6832 a_45124_376 VDD 0.259071f
C6833 a_47564_n7941 VDD 0.315469f
C6834 a_21940_n11684 a_23949_n12996 0.03954f
C6835 a_40620_n11077 VDD 0.343849f
C6836 a_32152_n13692 a_31960_n13648 0.934191f
C6837 a_32916_n15304 a_33004_n15348 0.285629f
C6838 a_23404_816 a_25524_n708 0.575323f
C6839 a_38380_n17349 VDD 0.342527f
C6840 a_34820_n16872 a_34908_n16916 0.285629f
C6841 a_31324_n16916 a_31772_n16916 0.013103f
C6842 a_24631_n3588 a_28144_n4708 0.263666f
C6843 a_42212_n20008 VDD 0.206217f
C6844 a_28492_332 a_29812_860 0.127939f
C6845 a_38733_n5431 a_39357_n5364 0.104193f
C6846 a_36773_n5468 a_37372_n5940 0.019402f
C6847 a_22444_n5156 a_26943_n7442 0.010531f
C6848 a_23479_n5156 a_24264_n6976 0.012448f
C6849 a_29123_n6679 a_31919_n9032 0.040884f
C6850 a_25612_n6679 a_33832_n8572 0.19454f
C6851 a_47028_n18820 a_47476_n18820 0.013276f
C6852 a_30584_n1954 VDD 0.611084f
C6853 a_46332_n20485 a_46244_n20388 0.285629f
C6854 a_46108_n9076 a_46556_n9076 0.012552f
C6855 a_47812_n9032 a_47900_n9076 0.285629f
C6856 a_39612_n4805 VDD 0.30038f
C6857 a_26531_n8639 VDD 0.318274f
C6858 a_40508_n12212 a_40956_n12212 0.012882f
C6859 a_46580_n10980 VDD 0.209016f
C6860 a_42604_n2020 a_45772_n101 0.021166f
C6861 a_36052_n14116 VDD 0.203482f
C6862 a_46020_n1572 a_46020_n2760 0.05841f
C6863 a_32432_n2689 a_32780_n2672 0.401636f
C6864 a_40420_n15304 a_40868_n15304 0.013276f
C6865 a_39188_n17252 VDD 0.211136f
C6866 a_38628_n16872 a_38268_n16916 0.087066f
C6867 a_42212_n4328 a_42660_n4328 0.013276f
C6868 a_30204_n20485 VDD 0.333707f
C6869 a_33533_908 a_30104_n1148 0.025895f
C6870 a_35119_398 a_35816_n174 0.212536f
C6871 a_35356_n18484 a_35804_n18484 0.012882f
C6872 a_29612_n8292 a_25612_n6679 0.088118f
C6873 a_26084_n20008 a_25724_n20052 0.087066f
C6874 a_28764_n8247 a_30228_n8203 0.487064f
C6875 a_43196_n7508 a_43084_n7941 0.026339f
C6876 a_34953_n1572 VDD 0.439779f
C6877 a_46244_n20388 a_46692_n20388 0.013276f
C6878 a_23564_n8292 a_24684_n16432 0.010489f
C6879 a_42660_n13736 CLK 0.017841f
C6880 a_42212_n9032 VDD 0.206217f
C6881 a_43196_n13780 a_43644_n13780 0.012882f
C6882 a_41092_n2760 a_40732_n2804 0.087174f
C6883 a_34796_n15348 a_34796_n15781 0.05841f
C6884 a_27628_n18484 VDD 0.329378f
C6885 a_45124_n16872 a_45572_n16872 0.013276f
C6886 a_39544_420 a_40260_n408 0.033597f
C6887 a_30564_n20388 VDD 0.208832f
C6888 a_42660_n18440 a_42300_n18484 0.087066f
C6889 a_23619_n6724 a_23949_n6724 0.538085f
C6890 a_32580_n20008 a_33028_n20008 0.013276f
C6891 a_31292_n2804 VDD 0.819314f
C6892 a_37820_n5940 VDD 0.331204f
C6893 a_25642_n9816 VDD 0.773325f
C6894 a_28121_n10980 a_28744_n14432 0.064531f
C6895 a_46916_n12168 VDD 0.205962f
C6896 a_26532_n14437 a_27192_n14286 0.096102f
C6897 a_39612_n13780 a_39724_n14213 0.026339f
C6898 a_46916_n1192 a_47364_n1192 0.013276f
C6899 a_45572_n1192 a_45660_n1236 0.285629f
C6900 a_39164_n15348 VDD 0.319301f
C6901 a_46916_n2760 a_46556_n2804 0.086742f
C6902 a_41852_n15348 a_41740_n15781 0.026339f
C6903 a_23036_n15781 a_22948_n15684 0.285629f
C6904 a_22052_1944 a_25084_1564 0.069988f
C6905 a_41764_n18440 VDD 0.206217f
C6906 a_24672_n11339 a_25237_n5895 0.257677f
C6907 a_44092_n16916 a_43980_n17349 0.026339f
C6908 a_39164_n4372 a_39164_n4805 0.05841f
C6909 a_23479_n5156 a_23207_n4708 0.022054f
C6910 a_47812_n18440 a_47900_n18484 0.285629f
C6911 a_46108_n18484 a_46556_n18484 0.012552f
C6912 a_37620_n7844 a_38068_n7844 0.013276f
C6913 a_44876_n7941 a_45236_n7844 0.087066f
C6914 a_42548_n10980 CLK 0.029747f
C6915 a_43420_n2804 VDD 0.317371f
C6916 a_38380_n9509 a_38740_n9412 0.087174f
C6917 a_21692_2431 VDD 1.36873f
C6918 a_29559_n6456 VDD 1.33811f
C6919 a_23564_n11428 a_24152_n11680 0.053516f
C6920 a_44876_n11077 a_45324_n11077 0.012882f
C6921 a_37036_n11077 a_37396_n10980 0.087174f
C6922 a_41740_n9509 VDD 0.313885f
C6923 a_35468_n12645 VDD 0.315889f
C6924 a_35692_n14213 a_36140_n14213 0.012882f
C6925 a_35244_n15781 VDD 0.296789f
C6926 a_42972_n2804 a_43084_n3237 0.026339f
C6927 a_25084_1564 a_26692_1564 0.010139f
C6928 a_26060_n18917 VDD 0.317718f
C6929 a_42636_n17349 a_43084_n17349 0.012882f
C6930 a_32108_n17349 a_32020_n17252 0.285629f
C6931 a_39412_n6276 a_39860_n6276 0.013276f
C6932 a_44876_n6373 a_44788_n6276 0.285629f
C6933 a_42660_n20008 a_42748_n20052 0.285629f
C6934 a_38716_n20052 a_39164_n20052 0.012882f
C6935 a_23479_n5156 a_26563_n12212 0.335147f
C6936 a_34552_n3140 VDD 0.360568f
C6937 a_32581_n9860 a_31872_n10529 0.050206f
C6938 a_41652_n9412 a_42100_n9412 0.013276f
C6939 a_26284_1564 VDD 0.010676f
C6940 a_45684_n6276 VDD 0.212747f
C6941 a_48012_n11077 a_47924_n10980 0.285629f
C6942 a_47924_n9412 VDD 0.21239f
C6943 a_42188_n12645 a_42548_n12548 0.087066f
C6944 a_39412_n12548 VDD 0.210723f
C6945 a_37932_n14213 a_38292_n14116 0.087066f
C6946 a_39636_n15684 VDD 0.209407f
C6947 a_33364_n15684 a_33812_n15684 0.013276f
C6948 a_28568_n16066 a_28548_n16872 0.014197f
C6949 a_42188_n15781 a_42100_n15684 0.285629f
C6950 a_29744_1564 a_30604_1515 0.882105f
C6951 a_47564_n18917 VDD 0.315469f
C6952 a_43980_n4805 a_44428_n4805 0.012882f
C6953 a_24672_n11339 a_24233_n5548 0.080017f
C6954 a_23228_n6679 a_22264_n5852 0.036868f
C6955 a_43084_n17349 a_43444_n17252 0.087066f
C6956 a_22052_n6980 a_24681_n7116 0.019043f
C6957 a_27852_n18917 a_28212_n18820 0.087066f
C6958 a_23324_n7420 a_23016_n7376 0.934191f
C6959 a_27988_n4328 a_27279_n12146 0.010988f
C6960 a_41292_n18917 a_41740_n18917 0.012882f
C6961 a_25860_n9032 a_25573_n12167 0.029991f
C6962 a_42748_n12212 CLK 0.012909f
C6963 a_46132_n3140 VDD 0.210512f
C6964 a_43416_1248 VDD 1.35109f
C6965 a_42660_n15304 CLK 0.017841f
C6966 a_37284_n7464 VDD 0.229013f
C6967 a_23564_n11428 a_21872_n12530 0.021744f
C6968 a_30808_n10600 VDD 0.608038f
C6969 a_28300_n15348 a_27852_n14990 0.122016f
C6970 a_40084_n14116 a_40532_n14116 0.013276f
C6971 a_34223_n1976 a_34953_n1572 0.212554f
C6972 a_33476_n16872 VDD 0.207033f
C6973 a_39412_n3140 a_39860_n3140 0.013276f
C6974 a_44428_n3237 a_44340_n3140 0.285629f
C6975 a_24631_n3588 a_26607_n3544 0.019779f
C6976 a_35849_n1192 a_36192_1248 0.10874f
C6977 a_42548_n18820 VDD 0.206098f
C6978 a_43444_n17252 a_43892_n17252 0.013276f
C6979 a_38828_n18917 a_38740_n18820 0.285629f
C6980 a_31799_n7508 a_32455_n7420 0.510371f
C6981 a_27055_n1192 VDD 0.575712f
C6982 a_34460_n20485 a_34908_n20485 0.013103f
C6983 a_33416_n4240 VDD 0.243199f
C6984 a_34271_376 VDD 0.694806f
C6985 a_47900_n7508 VDD 0.335152f
C6986 a_31279_n11728 a_30787_n12167 0.10971f
C6987 a_28927_n10160 a_30159_n13296 0.093895f
C6988 a_45660_n10644 VDD 0.320877f
C6989 a_27302_n13160 a_27526_n13714 0.75472f
C6990 a_38716_n13780 VDD 0.321613f
C6991 a_22948_n14820 a_23708_n15216 0.011851f
C6992 a_43332_n1572 a_43780_n1572 0.013276f
C6993 a_32860_n2020 a_32984_n2672 0.02305f
C6994 a_40508_n16916 VDD 0.313885f
C6995 a_37844_n15684 a_37732_n16872 0.026657f
C6996 a_21604_n3844 a_22364_n4240 0.011851f
C6997 a_22016_n4257 a_22876_n4284 0.882105f
C6998 a_27964_n20052 VDD 0.323654f
C6999 a_24292_n18440 a_23932_n18484 0.087174f
C7000 a_41652_n6276 CLK 0.016191f
C7001 a_36052_n18820 a_36500_n18820 0.013276f
C7002 a_38180_n7464 a_37820_n7508 0.087066f
C7003 a_22052_n18820 a_22052_n20008 0.05841f
C7004 a_42660_n9032 a_42300_n9076 0.087066f
C7005 a_34908_n20485 a_34820_n20388 0.285629f
C7006 a_26631_7 a_26527_51 0.277491f
C7007 a_38268_n9076 a_38716_n9076 0.012882f
C7008 a_47900_n4372 VDD 0.335152f
C7009 a_44540_332 VDD 0.34328f
C7010 a_47116_n7941 VDD 0.315469f
C7011 a_22600_n12124 a_21872_n12530 0.040755f
C7012 a_38180_n12168 a_38628_n12168 0.013276f
C7013 a_40172_n11077 VDD 0.315469f
C7014 a_31559_n13692 a_31960_n13648 0.882105f
C7015 a_35604_n15304 a_36052_n15304 0.013276f
C7016 a_25547_n2445 a_25139_n2704 0.056679f
C7017 a_31324_n4372 a_31348_n1931 0.216152f
C7018 a_37932_n17349 VDD 0.327654f
C7019 a_34820_n16872 a_34460_n16916 0.086905f
C7020 a_41764_n20008 VDD 0.206217f
C7021 a_22444_n5156 a_26719_n7464 0.010633f
C7022 a_32132_n18440 a_32580_n18440 0.013276f
C7023 a_23479_n5156 a_24681_n7116 0.02171f
C7024 a_29123_n6679 a_30900_n9032 0.74599f
C7025 a_44540_n7508 a_45124_n7464 0.016748f
C7026 a_29519_n1976 VDD 0.306953f
C7027 a_25831_n11428 a_34392_n9815 0.018612f
C7028 a_45884_n20485 a_46244_n20388 0.087174f
C7029 a_34820_n20388 a_35268_n20388 0.013276f
C7030 a_47812_n9032 a_47452_n9076 0.086635f
C7031 a_39164_n4805 VDD 0.302205f
C7032 a_42300_n10644 a_42748_n10644 0.012882f
C7033 a_23816_n8544 VDD 1.36785f
C7034 a_46132_n10980 VDD 0.210512f
C7035 a_45660_332 a_45772_n101 0.026339f
C7036 a_47197_908 a_47116_n101 0.029599f
C7037 a_39972_n13736 a_40420_n13736 0.013276f
C7038 a_35604_n14116 VDD 0.203482f
C7039 a_23608_n15260 a_24752_n16132 0.057444f
C7040 a_32860_n2020 a_22052_n4708 0.039953f
C7041 a_31392_n2760 a_32780_n2672 0.083829f
C7042 a_32432_n2689 a_33292_n2716 0.882105f
C7043 a_38740_n17252 VDD 0.213797f
C7044 a_41764_n16872 a_42212_n16872 0.013276f
C7045 a_33416_n4240 a_33868_n4240 0.026665f
C7046 a_38180_n16872 a_38268_n16916 0.285629f
C7047 a_29756_n20485 VDD 0.331916f
C7048 a_34895_376 a_35816_n174 0.01809f
C7049 a_32909_841 a_30104_n1148 0.02122f
C7050 a_42412_n5940 a_42860_n5940 0.013103f
C7051 a_21692_n20052 a_22140_n20052 0.012882f
C7052 a_25636_n20008 a_25724_n20052 0.285629f
C7053 a_42300_n9076 a_42188_n9509 0.026339f
C7054 a_22264_n10556 a_22220_n12996 0.820114f
C7055 a_42212_n13736 CLK 0.037136f
C7056 a_30871_n11728 a_28300_n15348 0.12801f
C7057 a_38268_n10644 a_38380_n11077 0.026339f
C7058 a_41764_n9032 VDD 0.206217f
C7059 a_38733_n727 a_39357_n660 0.104193f
C7060 a_24116_n15216 VDD 0.307009f
C7061 a_43196_n15348 a_43644_n15348 0.012882f
C7062 a_40644_n2760 a_40732_n2804 0.285629f
C7063 a_27180_n18484 VDD 0.333516f
C7064 a_44540_n4372 a_45124_n4328 0.016748f
C7065 a_38951_420 a_40260_n408 0.022815f
C7066 a_30116_n20388 VDD 0.206999f
C7067 a_38268_n18484 a_38716_n18484 0.012882f
C7068 a_42212_n18440 a_42300_n18484 0.285629f
C7069 a_37372_n5940 VDD 0.325054f
C7070 a_47452_n10644 a_47564_n11077 0.026339f
C7071 a_31961_n11340 a_31856_n11296 0.116059f
C7072 a_42948_n1976 a_43332_n1572 0.037522f
C7073 a_25237_n10599 VDD 0.502505f
C7074 a_46468_n12168 VDD 0.209055f
C7075 a_26532_n14437 a_26944_n14116 0.536965f
C7076 a_45572_n1192 a_45212_n1236 0.086905f
C7077 a_38716_n15348 VDD 0.321613f
C7078 a_46468_n2760 a_46556_n2804 0.285629f
C7079 a_22588_n15781 a_22948_n15684 0.086905f
C7080 a_41316_n18440 VDD 0.206217f
C7081 a_31212_n17349 a_31660_n17349 0.012222f
C7082 a_22444_n5156 a_22220_n9860 0.039352f
C7083 a_22544_n4690 a_23228_n6679 0.147748f
C7084 a_47924_376 a_48012_332 0.285629f
C7085 a_47812_n18440 a_47452_n18484 0.086635f
C7086 a_35356_n20052 a_35804_n20052 0.012882f
C7087 a_44876_n7941 a_44788_n7844 0.285629f
C7088 a_42100_n10980 CLK 0.020589f
C7089 a_42972_n2804 VDD 0.314361f
C7090 a_45772_n9509 a_46220_n9509 0.012882f
C7091 a_38380_n9509 a_38292_n9412 0.285629f
C7092 a_29211_n6724 VDD 0.47419f
C7093 a_37036_n11077 a_36948_n10980 0.285629f
C7094 a_24965_n9860 a_22016_n13665 0.053229f
C7095 a_41292_n9509 VDD 0.318502f
C7096 a_39500_n12645 a_39948_n12645 0.012222f
C7097 a_35020_n12645 VDD 0.327618f
C7098 a_25647_n1976 a_26271_n1400 0.104193f
C7099 a_34796_n15781 VDD 0.296789f
C7100 a_39276_n15781 a_39724_n15781 0.012882f
C7101 a_27337_n3140 a_25600_n5895 0.110889f
C7102 a_25612_n18917 VDD 0.325019f
C7103 a_31660_n17349 a_32020_n17252 0.086742f
C7104 a_24492_n5156 a_25573_n12167 0.186858f
C7105 a_44428_n6373 a_44788_n6276 0.087066f
C7106 a_30092_n18917 a_30540_n18917 0.012882f
C7107 a_42660_n20008 a_42300_n20052 0.087066f
C7108 a_34348_n3140 VDD 0.010384f
C7109 a_26796_1515 VDD 0.2446f
C7110 a_45236_n6276 VDD 0.229781f
C7111 a_47564_n11077 a_47924_n10980 0.087066f
C7112 a_39636_n10980 a_40084_n10980 0.013276f
C7113 a_29744_n10980 a_30787_n12167 0.012356f
C7114 a_47476_n9412 VDD 0.206217f
C7115 a_42188_n12645 a_42100_n12548 0.285629f
C7116 a_38964_n12548 VDD 0.212805f
C7117 a_37932_n14213 a_37844_n14116 0.285629f
C7118 a_46220_n14213 a_46668_n14213 0.012882f
C7119 a_39188_n15684 VDD 0.211136f
C7120 a_41740_n15781 a_42100_n15684 0.087066f
C7121 a_29332_1243 a_30296_1564 0.08126f
C7122 a_29744_1564 a_28836_376 0.391901f
C7123 a_47116_n18917 VDD 0.315469f
C7124 a_32020_n17252 a_32468_n17252 0.013276f
C7125 a_43084_n17349 a_42996_n17252 0.285629f
C7126 a_24492_n5156 a_23816_n5408 0.037526f
C7127 a_23228_n6679 a_22016_n5825 0.024424f
C7128 a_22544_n4690 a_22772_n5808 0.019536f
C7129 a_27852_n18917 a_27764_n18820 0.285629f
C7130 a_47812_n20008 a_47900_n20052 0.285629f
C7131 a_46108_n20052 a_46556_n20052 0.012552f
C7132 a_42100_n7844 a_42212_n9032 0.026657f
C7133 a_42300_n12212 CLK 0.048577f
C7134 a_45684_n3140 VDD 0.212747f
C7135 a_22876_n10556 a_22772_n10512 0.026665f
C7136 a_23564_n8292 a_23949_n12996 0.028852f
C7137 a_42372_1564 VDD 0.298894f
C7138 a_42212_n15304 CLK 0.037136f
C7139 a_22352_n12097 a_24152_n11680 0.510371f
C7140 a_23564_n11428 a_23619_n12996 0.047156f
C7141 a_43892_n12548 a_44340_n12548 0.013276f
C7142 a_28300_n15348 a_27404_n14990 0.307662f
C7143 a_30555_n13780 VDD 0.493833f
C7144 a_33999_n1400 a_34953_n1572 0.014822f
C7145 a_22052_1944 OUT[0] 0.265324f
C7146 a_33028_n16872 VDD 0.212051f
C7147 a_43892_n15684 a_44340_n15684 0.013276f
C7148 a_43980_n3237 a_44340_n3140 0.087066f
C7149 a_24631_n3588 a_26383_n2968 0.013293f
C7150 a_22096_376 a_22340_376 0.014807f
C7151 a_42100_n18820 VDD 0.206098f
C7152 a_42548_n4708 a_42996_n4708 0.013276f
C7153 a_31799_n7508 a_32560_n7020 0.042802f
C7154 a_38380_n18917 a_38740_n18820 0.087066f
C7155 a_31451_n7508 a_32455_n7420 0.020455f
C7156 a_32262_n452 VDD 0.656973f
C7157 a_29123_n6679 a_29176_n7819 0.010396f
C7158 a_26431_n1192 VDD 0.714427f
C7159 a_44509_n452 a_42948_n1976 0.465348f
C7160 a_28225_n4327 VDD 0.966776f
C7161 a_32581_n9860 a_31961_n11340 0.019421f
C7162 a_30808_n10116 a_31872_n10529 0.351723f
C7163 a_31460_n10116 a_32424_n10512 0.08126f
C7164 a_34403_332 VDD 0.554918f
C7165 a_47452_n7508 VDD 0.313885f
C7166 a_44340_n10980 a_44452_n12168 0.026657f
C7167 a_45212_n10644 VDD 0.342281f
C7168 a_38268_n13780 VDD 0.356784f
C7169 a_22948_n14820 a_24220_n15260 0.05539f
C7170 a_32860_n2020 a_32780_n2672 0.018082f
C7171 a_40060_n16916 VDD 0.314419f
C7172 a_22016_n4257 a_21792_n7464 0.369876f
C7173 a_21604_n3844 a_22876_n4284 0.05539f
C7174 a_27516_n20052 VDD 0.316938f
C7175 a_40420_n4708 a_40532_n5896 0.026657f
C7176 a_27540_n18440 a_27988_n18440 0.013276f
C7177 a_23844_n18440 a_23932_n18484 0.285629f
C7178 a_41204_n6276 CLK 0.015237f
C7179 a_41316_n7464 a_41764_n7464 0.013276f
C7180 a_37732_n7464 a_37820_n7508 0.285629f
C7181 a_26631_7 a_27224_n62 0.361958f
C7182 a_42212_n9032 a_42300_n9076 0.285629f
C7183 a_45436_n20485 a_45884_n20485 0.013103f
C7184 a_34460_n20485 a_34820_n20388 0.087174f
C7185 a_47452_n4372 VDD 0.313885f
C7186 a_39076_n10600 a_39524_n10600 0.013276f
C7187 a_46668_n7941 VDD 0.318039f
C7188 a_39724_n11077 VDD 0.318714f
C7189 a_31664_n13292 a_31960_n13648 0.05539f
C7190 a_31459_n14564 VDD 0.35969f
C7191 a_24771_n2804 a_25139_n2704 0.569174f
C7192 a_23507_n2759 a_23319_n2759 0.255962f
C7193 a_31324_n4372 a_27988_n4328 0.035234f
C7194 a_37484_n17349 VDD 0.322148f
C7195 a_34372_n16872 a_34460_n16916 0.285629f
C7196 a_30876_n16916 a_31324_n16916 0.013103f
C7197 a_22052_n4708 a_23887_n5156 0.013478f
C7198 a_41316_n20008 VDD 0.206217f
C7199 a_22444_n5156 a_26095_n7464 0.012149f
C7200 a_38403_n5503 a_38733_n5431 0.538085f
C7201 a_46580_n18820 a_47028_n18820 0.013276f
C7202 a_22220_n9860 a_21604_n10116 0.036078f
C7203 a_23479_n5156 a_27485_n10068 0.030453f
C7204 a_24672_n11339 a_23816_n10112 0.024322f
C7205 a_29295_n1400 VDD 0.574776f
C7206 a_45660_n9076 a_46108_n9076 0.012552f
C7207 a_45884_n20485 a_45796_n20388 0.285629f
C7208 a_25831_n11428 a_33494_n9860 0.025562f
C7209 a_47364_n9032 a_47452_n9076 0.285629f
C7210 a_38716_n4805 VDD 0.335795f
C7211 a_24233_n8684 VDD 0.498506f
C7212 a_44452_n12168 a_44540_n12212 0.285629f
C7213 a_40060_n12212 a_40508_n12212 0.012882f
C7214 a_31279_n11728 a_31459_n12996 0.21401f
C7215 a_45684_n10980 VDD 0.212747f
C7216 a_42604_n2020 a_42948_n1976 0.177017f
C7217 a_30104_n1148 a_30781_n452 0.016705f
C7218 a_35156_n14116 VDD 0.203482f
C7219 a_39972_n15304 a_40420_n15304 0.013276f
C7220 a_45572_n1572 a_45572_n2760 0.05841f
C7221 a_38292_n17252 VDD 0.243749f
C7222 a_41764_n4328 a_42212_n4328 0.013276f
C7223 a_38180_n16872 a_37820_n16916 0.087066f
C7224 a_28636_n16916 a_28524_n17349 0.026339f
C7225 a_32579_769 a_30104_n1148 0.019285f
C7226 a_29308_n20485 VDD 0.335406f
C7227 a_34908_n18484 a_35356_n18484 0.012882f
C7228 a_26631_7 VDD 0.805322f
C7229 a_25636_n20008 a_25276_n20052 0.087066f
C7230 a_42748_n7508 a_42636_n7941 0.026339f
C7231 a_32100_n1976 VDD 0.830948f
C7232 a_43555_n452 a_42948_n1976 0.034477f
C7233 a_45796_n20388 a_46244_n20388 0.013276f
C7234 a_24965_n9860 a_25831_n12996 0.02806f
C7235 a_41316_n9032 VDD 0.206217f
C7236 a_42748_n13780 a_43196_n13780 0.012882f
C7237 a_25472_n14816 VDD 0.023744f
C7238 a_34348_n15348 a_34348_n15781 0.05841f
C7239 a_43780_n2760 a_44228_n2760 0.013276f
C7240 a_26172_n18484 VDD 0.332466f
C7241 a_36700_n16916 a_36588_n17349 0.026339f
C7242 a_44540_n16916 a_45124_n16872 0.016748f
C7243 a_27988_n20388 a_27852_n18917 0.027118f
C7244 a_29668_n20388 VDD 0.204779f
C7245 a_39056_820 a_40260_n408 0.021298f
C7246 a_42212_n18440 a_41852_n18484 0.087066f
C7247 a_42636_n7941 CLK 0.01698f
C7248 a_32132_n20008 a_32580_n20008 0.013276f
C7249 a_32189_n9860 a_32581_n9860 0.466799f
C7250 a_44116_n5896 VDD 0.2198f
C7251 a_31544_n11296 a_31856_n11296 0.119687f
C7252 a_24965_n9860 VDD 0.876106f
C7253 a_28040_n12493 a_28492_n12548 0.026665f
C7254 a_46020_n12168 VDD 0.210736f
C7255 a_46468_n1192 a_46916_n1192 0.013276f
C7256 a_39164_n13780 a_39276_n14213 0.026339f
C7257 a_45124_n1192 a_45212_n1236 0.285629f
C7258 a_38268_n15348 VDD 0.356784f
C7259 a_46468_n2760 a_46108_n2804 0.086905f
C7260 a_41404_n15348 a_41292_n15781 0.026339f
C7261 a_22588_n15781 a_22500_n15684 0.285629f
C7262 a_40652_n1572 a_45572_n1572 0.038441f
C7263 a_21692_2431 a_25084_1564 1.94336f
C7264 a_40868_n18440 VDD 0.208618f
C7265 a_43644_n16916 a_43532_n17349 0.026339f
C7266 a_47364_n18440 a_47452_n18484 0.285629f
C7267 a_45660_n18484 a_46108_n18484 0.012552f
C7268 a_44428_n7941 a_44788_n7844 0.087066f
C7269 a_37172_n7844 a_37620_n7844 0.013276f
C7270 a_25972_n6276 a_25020_n11383 0.010178f
C7271 a_42524_n2804 VDD 0.314361f
C7272 a_25860_n9032 a_24964_n14116 0.014739f
C7273 a_37932_n9509 a_38292_n9412 0.087174f
C7274 a_25573_n12167 a_23564_n11428 0.829302f
C7275 a_36588_n11077 a_36948_n10980 0.087174f
C7276 a_24965_n9860 a_21604_n13252 0.010201f
C7277 a_44428_n11077 a_44876_n11077 0.012882f
C7278 a_40620_n9509 VDD 0.344269f
C7279 a_34572_n12645 VDD 0.316938f
C7280 a_35244_n14213 a_35692_n14213 0.012882f
C7281 a_34348_n15781 VDD 0.296789f
C7282 a_22820_n2804 a_33015_n4284 0.047274f
C7283 a_42524_n2804 a_42636_n3237 0.026339f
C7284 a_24631_n3588 a_22164_n2760 0.194717f
C7285 a_28736_1944 a_28153_1204 0.031565f
C7286 a_24828_n18917 VDD 0.337122f
C7287 a_42188_n17349 a_42636_n17349 0.012882f
C7288 a_47900_n4372 a_48012_n4805 0.026339f
C7289 a_31660_n17349 a_31572_n17252 0.285629f
C7290 a_24672_n11339 a_25860_n9032 0.010665f
C7291 a_44428_n6373 a_44340_n6276 0.285629f
C7292 a_25612_n6679 a_30036_n7464 0.022442f
C7293 a_38268_n20052 a_38716_n20052 0.012882f
C7294 a_42212_n20008 a_42300_n20052 0.285629f
C7295 a_34860_n3189 VDD 0.243199f
C7296 a_32581_n9860 a_30808_n10116 0.024997f
C7297 a_22096_376 VDD 0.283746f
C7298 a_41204_n9412 a_41652_n9412 0.013276f
C7299 a_44788_n6276 VDD 0.22479f
C7300 a_27281_n16854 a_27820_n16432 0.241389f
C7301 a_28927_n10160 a_33488_n12996 0.565925f
C7302 a_47564_n11077 a_47476_n10980 0.285629f
C7303 a_47028_n9412 VDD 0.206217f
C7304 a_41740_n12645 a_42100_n12548 0.087066f
C7305 a_38516_n12548 VDD 0.216736f
C7306 a_37484_n14213 a_37844_n14116 0.087066f
C7307 a_38740_n15684 VDD 0.213797f
C7308 a_43644_n705 OUT[5] 0.012713f
C7309 a_41740_n15781 a_41652_n15684 0.285629f
C7310 a_29332_1243 a_30092_1564 0.011851f
C7311 a_46668_n18917 VDD 0.318039f
C7312 a_23887_n5156 a_23816_n5408 0.061392f
C7313 a_42636_n17349 a_42996_n17252 0.087066f
C7314 a_43532_n4805 a_43980_n4805 0.012882f
C7315 a_24492_n5156 a_24233_n5548 0.038689f
C7316 a_23228_n6679 a_21604_n5412 0.031222f
C7317 a_22712_n7420 a_22812_n7376 0.092119f
C7318 a_22464_n7393 a_23016_n7376 0.361958f
C7319 a_27404_n18917 a_27764_n18820 0.087066f
C7320 a_47812_n20008 a_47452_n20052 0.086635f
C7321 a_41852_n12212 CLK 0.013107f
C7322 a_45236_n3140 VDD 0.229781f
C7323 a_42168_1564 VDD 0.360568f
C7324 a_34176_n6976 VDD 0.010384f
C7325 a_28300_n15348 a_31760_n12168 0.500353f
C7326 a_22352_n12097 a_24569_n11820 0.020455f
C7327 a_21940_n11684 a_24152_n11680 0.042802f
C7328 a_22700_n12080 a_22904_n12080 0.048436f
C7329 a_33984_n10112 VDD 0.022335f
C7330 a_30159_n13296 VDD 1.13498f
C7331 a_28752_n15348 a_28212_n15303 0.010551f
C7332 a_39636_n14116 a_40084_n14116 0.013276f
C7333 a_32580_n16872 VDD 0.213022f
C7334 a_43980_n3237 a_43892_n3140 0.285629f
C7335 a_37396_1205 a_37844_1564 0.21055f
C7336 a_25524_1243 a_25817_804 0.04091f
C7337 a_41652_n18820 VDD 0.206098f
C7338 a_42996_n17252 a_43444_n17252 0.013276f
C7339 a_23479_n5156 a_27526_n9816 0.018948f
C7340 a_31451_n7508 a_32560_n7020 0.019043f
C7341 a_38380_n18917 a_38292_n18820 0.285629f
C7342 a_27988_n20388 XRST 0.058012f
C7343 a_34012_n20485 a_34460_n20485 0.013103f
C7344 a_43885_n452 a_42948_n1976 0.088306f
C7345 a_32911_n4240 VDD 0.022892f
C7346 a_31460_n10116 a_32220_n10512 0.011851f
C7347 a_32581_n9860 a_31544_n11296 0.035551f
C7348 a_33533_908 VDD 0.705267f
C7349 a_47004_n7508 VDD 0.313885f
C7350 a_43644_n705 a_42948_n1976 0.206043f
C7351 a_47812_n10600 VDD 0.211703f
C7352 a_25831_n12996 a_25636_n14520 0.057189f
C7353 a_26470_n13736 a_27302_n13160 0.106585f
C7354 a_37820_n13780 VDD 0.322978f
C7355 a_22948_n14820 a_23608_n15260 0.113808f
C7356 a_39612_n16916 VDD 0.317476f
C7357 a_28548_n16872 a_28636_n16916 0.285629f
C7358 a_37396_n15684 a_37284_n16872 0.026657f
C7359 a_21604_n3844 a_21792_n7464 0.109028f
C7360 a_27068_n20052 VDD 0.328902f
C7361 a_23844_n18440 a_23484_n18484 0.087174f
C7362 a_22016_n5825 a_24128_n5408 0.277491f
C7363 a_27988_n4328 a_27281_n16854 0.040235f
C7364 a_40308_n6276 CLK 0.014457f
C7365 a_21604_n18820 a_21604_n20008 0.05841f
C7366 a_37732_n7464 a_37372_n7508 0.087066f
C7367 a_35604_n18820 a_36052_n18820 0.013276f
C7368 a_34460_n20485 a_34372_n20388 0.285629f
C7369 a_26736_n364 a_27224_n62 0.08126f
C7370 a_42212_n9032 a_41852_n9076 0.087066f
C7371 a_37820_n9076 a_38268_n9076 0.012882f
C7372 a_23564_n8292 a_24128_n10112 0.049334f
C7373 a_25975_n184 a_26527_51 0.119687f
C7374 a_47004_n4372 VDD 0.313885f
C7375 a_39804_464 VDD 0.299466f
C7376 a_46220_n7941 VDD 0.31977f
C7377 a_22600_n12124 a_21772_n12996 0.473936f
C7378 a_37732_n12168 a_38180_n12168 0.013276f
C7379 a_42636_n18917 CLK 0.01698f
C7380 a_39276_n11077 VDD 0.320362f
C7381 a_31559_n13692 a_31455_n13648 0.277491f
C7382 a_25636_n14520 VDD 0.833044f
C7383 a_37221_n3543 a_37452_n3888 0.075587f
C7384 a_35156_n15304 a_35604_n15304 0.013276f
C7385 a_34248_n3310 a_34232_n2272 0.055219f
C7386 a_27316_n14820 a_28212_n15303 0.01161f
C7387 a_37036_n17349 VDD 0.334604f
C7388 a_22052_n4708 a_23479_n5156 0.010602f
C7389 a_34372_n16872 a_34012_n16916 0.086905f
C7390 a_40868_n20008 VDD 0.208618f
C7391 a_31684_n18440 a_32132_n18440 0.013276f
C7392 a_44340_n17252 a_44452_n18440 0.026657f
C7393 a_47924_n4708 a_47812_n5896 0.026657f
C7394 a_23887_n5156 a_23016_n7376 0.031986f
C7395 a_24672_n11339 a_22712_n7420 0.028662f
C7396 a_24672_n11339 a_24233_n10252 0.045757f
C7397 a_23479_n5156 a_26861_n10135 0.069029f
C7398 a_44092_n7508 a_44540_n7508 0.012001f
C7399 a_25972_n6276 a_32767_n9010 0.020458f
C7400 a_47364_n9032 a_47004_n9076 0.086742f
C7401 a_45436_n20485 a_45796_n20388 0.087174f
C7402 a_34372_n20388 a_34820_n20388 0.013276f
C7403 a_38268_n4805 VDD 0.371393f
C7404 a_41852_n10644 a_42300_n10644 0.012882f
C7405 a_44452_n12168 a_44092_n12212 0.086635f
C7406 a_28009_n12168 a_29360_n12864 0.114166f
C7407 a_45236_n10980 VDD 0.229781f
C7408 a_27526_n13714 a_26532_n14437 0.031746f
C7409 a_46573_841 a_46668_n101 0.025027f
C7410 a_45212_332 a_45324_n101 0.026339f
C7411 a_39524_n13736 a_39972_n13736 0.013276f
C7412 a_34708_n14116 VDD 0.203482f
C7413 a_32020_n2276 a_34232_n2272 0.042803f
C7414 a_31392_n2760 a_32432_n2689 0.348372f
C7415 a_40652_n1572 a_45660_n1236 0.022582f
C7416 a_37844_n17252 VDD 0.214349f
C7417 a_23564_n20836 a_24292_n18440 0.017841f
C7418 a_41316_n16872 a_41764_n16872 0.013276f
C7419 a_37732_n16872 a_37820_n16916 0.285629f
C7420 a_28300_n20485 VDD 0.333555f
C7421 a_41964_n5940 a_42412_n5940 0.013103f
C7422 a_25188_n20008 a_25276_n20052 0.285629f
C7423 a_27597_n8292 a_28764_n8247 0.010748f
C7424 a_26736_n364 VDD 1.7793f
C7425 a_42860_n101 a_42948_n1976 0.022318f
C7426 a_41852_n9076 a_41740_n9509 0.026339f
C7427 a_47924_n4708 VDD 0.21239f
C7428 a_37820_n10644 a_37932_n11077 0.026339f
C7429 a_24760_n11383 a_24964_n14116 0.014899f
C7430 a_21772_n9860 a_21892_n12952 0.027496f
C7431 a_40868_n9032 VDD 0.208618f
C7432 a_47452_n12212 a_47900_n12212 0.012001f
C7433 a_29920_n12168 VDD 0.010055f
C7434 a_38403_n799 a_38733_n727 0.538085f
C7435 a_39308_n452 a_41533_n727 0.024548f
C7436 a_42748_n15348 a_43196_n15348 0.012882f
C7437 a_31324_n4372 a_32020_n2276 0.01069f
C7438 a_25724_n18484 VDD 0.320117f
C7439 a_44092_n4372 a_44540_n4372 0.012001f
C7440 a_27988_n20388 a_27404_n18917 0.030758f
C7441 a_29220_n20388 VDD 0.225668f
C7442 a_40196_1944 OUT[4] 0.225001f
C7443 a_24492_n5156 a_28764_n8247 0.014373f
C7444 a_37820_n18484 a_38268_n18484 0.012882f
C7445 a_41764_n18440 a_41852_n18484 0.285629f
C7446 a_42188_n7941 CLK 0.050454f
C7447 a_23479_n5156 a_26543_n11384 0.021753f
C7448 a_24672_n11339 a_24760_n11383 0.251198f
C7449 a_39948_n7941 a_40396_n7941 0.012222f
C7450 a_27348_n2672 VDD 0.01368f
C7451 a_31565_n9860 a_32581_n9860 0.059672f
C7452 a_43668_n5896 VDD 0.212309f
C7453 a_47004_n10644 a_47116_n11077 0.026339f
C7454 a_31544_n11296 a_31961_n11340 0.633318f
C7455 a_24573_n9860 VDD 0.837993f
C7456 a_27744_n12908 a_29360_n12864 0.011851f
C7457 a_45572_n12168 VDD 0.213324f
C7458 a_37820_n15348 VDD 0.322978f
C7459 a_22140_n15781 a_22500_n15684 0.086905f
C7460 a_46020_n2760 a_46108_n2804 0.285629f
C7461 a_47364_n2760 a_47812_n2760 0.013276f
C7462 a_42604_n2020 a_46468_n1192 0.017841f
C7463 a_40652_n1572 a_45124_n1572 0.021187f
C7464 a_40420_n18440 VDD 0.205948f
C7465 a_30764_n17349 a_31212_n17349 0.013103f
C7466 a_24492_n5156 a_24672_n11339 0.026236f
C7467 a_22444_n5156 a_23228_n6679 0.013066f
C7468 a_47364_n18440 a_47004_n18484 0.086742f
C7469 a_44428_n7941 a_44340_n7844 0.285629f
C7470 a_34908_n20052 a_35356_n20052 0.012882f
C7471 a_42076_n2804 VDD 0.314361f
C7472 a_37932_n9509 a_37844_n9412 0.285629f
C7473 a_45324_n9509 a_45772_n9509 0.012882f
C7474 a_25972_n6276 VDD 1.32364f
C7475 a_40172_n9509 VDD 0.315889f
C7476 a_39052_n12645 a_39500_n12645 0.012222f
C7477 a_34124_n12645 VDD 0.311881f
C7478 a_27820_n16432 a_27988_n20388 0.691737f
C7479 a_33900_n15781 VDD 0.296789f
C7480 a_27672_n3543 a_28583_n3140 0.015754f
C7481 a_38828_n15781 a_39276_n15781 0.012882f
C7482 a_22820_n2804 a_33120_n3884 0.017389f
C7483 a_24380_n18917 VDD 0.315637f
C7484 a_22500_n1976 a_28153_1204 0.039552f
C7485 a_28736_1944 a_27736_1248 0.038332f
C7486 a_31212_n17349 a_31572_n17252 0.086742f
C7487 a_43980_n6373 a_44340_n6276 0.087066f
C7488 a_29644_n18917 a_30092_n18917 0.012882f
C7489 a_23479_n5156 a_25573_n12167 0.375631f
C7490 a_42212_n20008 a_41852_n20052 0.087066f
C7491 a_34000_n3140 VDD 0.797914f
C7492 a_39556_n4 a_39760_n4 0.033243f
C7493 a_25936_1564 VDD 0.806659f
C7494 a_44340_n6276 VDD 0.212126f
C7495 a_47116_n11077 a_47476_n10980 0.087066f
C7496 a_28927_n10160 a_32413_n12996 0.475806f
C7497 a_39188_n10980 a_39636_n10980 0.013276f
C7498 a_46580_n9412 VDD 0.209016f
C7499 a_41740_n12645 a_41652_n12548 0.285629f
C7500 a_38068_n12548 VDD 0.230258f
C7501 a_45772_n14213 a_46220_n14213 0.012882f
C7502 a_37484_n14213 a_37396_n14116 0.285629f
C7503 a_38292_n15684 VDD 0.243749f
C7504 a_41292_n15781 a_41652_n15684 0.087066f
C7505 a_40196_1944 a_41204_1243 0.095846f
C7506 a_29332_1243 a_30604_1515 0.05539f
C7507 a_46220_n18917 VDD 0.31977f
C7508 a_31572_n17252 a_32020_n17252 0.013276f
C7509 a_42636_n17349 a_42548_n17252 0.285629f
C7510 a_27404_n18917 a_27316_n18820 0.285629f
C7511 a_22464_n7393 a_22812_n7376 0.401636f
C7512 a_22052_n6980 a_23016_n7376 0.08126f
C7513 OUT[5] EOC 0.016184f
C7514 a_45660_n20052 a_46108_n20052 0.012552f
C7515 a_47364_n20008 a_47452_n20052 0.285629f
C7516 a_41652_n7844 a_41764_n9032 0.026657f
C7517 a_44788_n3140 VDD 0.22479f
C7518 a_25020_n11383 a_30871_n11728 0.355014f
C7519 a_24233_n10252 a_23816_n10112 0.633318f
C7520 a_22016_n10529 a_24128_n10112 0.277491f
C7521 a_41964_1564 VDD 0.010384f
C7522 a_21940_n11684 a_24569_n11820 0.019043f
C7523 a_23212_n12124 a_22904_n12080 0.934191f
C7524 a_43444_n12548 a_43892_n12548 0.013276f
C7525 a_32308_n1976 a_34248_n3310 0.038089f
C7526 a_24315_n2759 a_23319_n2759 0.064779f
C7527 a_41684_n1976 a_42244_n1572 0.302602f
C7528 a_32132_n16872 VDD 0.213947f
C7529 a_43444_n15684 a_43892_n15684 0.013276f
C7530 a_23564_n17700 a_23932_n16916 0.032404f
C7531 a_43532_n3237 a_43892_n3140 0.087066f
C7532 a_41204_n18820 VDD 0.226851f
C7533 a_42100_n4708 a_42548_n4708 0.013276f
C7534 a_37932_n18917 a_38292_n18820 0.087066f
C7535 a_24292_n18820 a_24740_n18820 0.013276f
C7536 a_25972_n6276 a_30676_n7844 0.714881f
C7537 a_23479_n5156 a_27302_n9816 0.083519f
C7538 a_31405_n452 VDD 0.770376f
C7539 a_23816_n704 VDD 1.36367f
C7540 a_43885_n452 a_44509_n452 0.104193f
C7541 a_33608_n4284 VDD 0.360568f
C7542 a_31460_n10116 a_32732_n10556 0.05539f
C7543 a_32909_841 VDD 0.594208f
C7544 a_46556_n7508 VDD 0.31705f
C7545 a_43892_n10980 a_44004_n12168 0.026657f
C7546 a_33686_n11592 a_33910_n12146 0.75472f
C7547 a_47364_n10600 VDD 0.205948f
C7548 a_43644_n705 a_44509_n452 0.013628f
C7549 a_23816_n13248 a_24128_n13248 0.119687f
C7550 a_37372_n13780 VDD 0.325523f
C7551 a_21692_n15348 a_22140_n15348 0.012222f
C7552 a_22948_n14820 a_23360_n15233 0.536965f
C7553 a_32860_n2020 a_32432_n2689 0.046548f
C7554 a_39164_n16916 VDD 0.319301f
C7555 a_21604_n3844 a_22016_n4257 0.536965f
C7556 a_43644_n705 a_45012_1564 0.274319f
C7557 a_33467_1116 a_33533_908 0.017118f
C7558 a_26620_n20052 VDD 0.328902f
C7559 a_22876_n5852 a_23816_n5408 0.056721f
C7560 a_23396_n18440 a_23484_n18484 0.285629f
C7561 a_39972_n4708 a_40084_n5896 0.026657f
C7562 a_27092_n18440 a_27540_n18440 0.013276f
C7563 a_39860_n6276 CLK 0.014484f
C7564 a_37284_n7464 a_37372_n7508 0.285629f
C7565 a_40868_n7464 a_41316_n7464 0.013276f
C7566 a_42548_n9412 CLK 0.029747f
C7567 a_44988_n20485 a_45436_n20485 0.013103f
C7568 a_34012_n20485 a_34372_n20388 0.087174f
C7569 a_41764_n9032 a_41852_n9076 0.285629f
C7570 a_25627_n452 a_26527_51 0.116059f
C7571 a_22264_n8988 a_22220_n12996 0.286379f
C7572 a_46556_n4372 VDD 0.31705f
C7573 a_38628_n10600 a_39076_n10600 0.013276f
C7574 a_23816_n10112 a_24760_n11383 0.027122f
C7575 a_45772_n7941 VDD 0.321879f
C7576 a_21940_n11684 a_23619_n12996 0.030938f
C7577 a_38828_n11077 VDD 0.322604f
C7578 a_42188_n18917 CLK 0.047331f
C7579 a_30903_n13780 a_31960_n13648 0.056721f
C7580 a_31559_n13692 a_32152_n13692 0.361958f
C7581 a_29056_n14432 VDD 0.022335f
C7582 a_24771_n2804 a_25547_n2445 0.153996f
C7583 a_23507_n2759 a_25139_n2704 0.021458f
C7584 a_34248_n3310 a_34649_n2412 0.058671f
C7585 a_36588_n17349 VDD 0.316762f
C7586 a_30428_n16916 a_30876_n16916 0.013103f
C7587 a_33924_n16872 a_34012_n16916 0.285629f
C7588 a_40420_n20008 VDD 0.205948f
C7589 a_45236_n4 a_45684_n4 0.013276f
C7590 a_23479_n5156 a_23016_n7376 0.010191f
C7591 a_25972_n6276 a_32543_n9032 0.029586f
C7592 a_46132_n18820 a_46580_n18820 0.013276f
C7593 a_23479_n5156 a_26531_n10207 0.02061f
C7594 a_27706_n1572 VDD 0.014238f
C7595 a_45212_n9076 a_45660_n9076 0.012552f
C7596 a_45436_n20485 a_45348_n20388 0.285629f
C7597 a_46916_n9032 a_47004_n9076 0.285629f
C7598 a_25831_n11428 a_32189_n9860 0.026608f
C7599 a_44004_n12168 a_44092_n12212 0.285629f
C7600 a_27281_n16854 a_27316_n14820 0.065239f
C7601 a_39612_n12212 a_40060_n12212 0.012882f
C7602 a_44788_n10980 VDD 0.22479f
C7603 a_27302_n13160 a_26532_n14437 0.04208f
C7604 a_30104_n1148 a_30451_n452 0.054397f
C7605 a_34260_n14116 VDD 0.203482f
C7606 a_39524_n15304 a_39972_n15304 0.013276f
C7607 a_45124_n1572 a_45124_n2760 0.05841f
C7608 a_32020_n2276 a_34649_n2412 0.019033f
C7609 a_40652_n1572 a_45212_n1236 0.029702f
C7610 a_37396_n17252 VDD 0.211702f
C7611 a_37732_n16872 a_37372_n16916 0.087066f
C7612 a_41316_n4328 a_41764_n4328 0.013276f
C7613 a_23564_n20836 a_23844_n18440 0.036527f
C7614 a_33608_n4284 a_33868_n4240 0.66083f
C7615 a_27540_n20747 VDD 0.463305f
C7616 a_43644_n705 a_42604_n2020 0.030792f
C7617 a_24631_n3588 a_30104_n1148 0.05018f
C7618 a_34460_n18484 a_34908_n18484 0.012882f
C7619 a_25975_n184 VDD 1.34345f
C7620 a_42300_n7508 a_42188_n7941 0.026339f
C7621 a_25188_n20008 a_24828_n20052 0.087066f
C7622 a_22712_n7420 a_25860_n9032 0.102125f
C7623 a_47900_n1669 VDD 0.318055f
C7624 a_45348_n20388 a_45796_n20388 0.013276f
C7625 a_43555_n452 a_43885_n452 0.538085f
C7626 a_21772_n9860 a_22220_n12996 0.032585f
C7627 a_47476_n4708 VDD 0.206217f
C7628 a_22264_n8988 a_22568_n13648 0.049352f
C7629 a_42660_n16872 CLK 0.017841f
C7630 a_40420_n9032 VDD 0.206217f
C7631 a_30599_n12167 VDD 1.01111f
C7632 a_43644_n705 a_43555_n452 0.054785f
C7633 a_42300_n13780 a_42748_n13780 0.012882f
C7634 a_27224_n62 a_27032_51 0.934191f
C7635 a_27852_n14990 VDD 0.61975f
C7636 a_39308_n452 a_41203_n799 0.239811f
C7637 a_38996_n408 a_39357_n660 0.034982f
C7638 a_33900_n15348 a_33900_n15781 0.05841f
C7639 a_23507_n2759 a_25600_n5895 0.153739f
C7640 a_43332_n2760 a_43780_n2760 0.013276f
C7641 a_31324_n4372 a_31292_n2804 0.576967f
C7642 a_25276_n18484 VDD 0.337006f
C7643 a_44092_n16916 a_44540_n16916 0.012001f
C7644 a_22052_n4708 a_22264_n5852 0.011359f
C7645 a_36252_n16916 a_36140_n17349 0.026339f
C7646 a_28212_n20388 VDD 0.126945f
C7647 a_41764_n18440 a_41404_n18484 0.087066f
C7648 a_41740_n7941 CLK 0.01075f
C7649 a_24672_n11339 a_23564_n11428 0.021115f
C7650 a_23479_n5156 a_26547_n12951 0.098988f
C7651 a_31684_n20008 a_32132_n20008 0.013276f
C7652 a_29992_n11150 a_32581_n9860 0.028587f
C7653 a_31565_n9860 a_32189_n9860 0.104193f
C7654 a_43220_n5896 VDD 0.209811f
C7655 a_28927_n10160 a_31760_n12168 0.374556f
C7656 a_23949_n9860 VDD 0.594438f
C7657 a_27744_n12908 a_30340_n12548 0.094068f
C7658 a_28232_n12606 a_28492_n12548 0.66083f
C7659 a_45124_n12168 VDD 0.26277f
C7660 a_38716_n13780 a_38828_n14213 0.026339f
C7661 a_46020_n1192 a_46468_n1192 0.013276f
C7662 a_37372_n15348 VDD 0.325523f
C7663 a_22140_n15781 a_22052_n15684 0.285629f
C7664 a_46020_n2760 a_45660_n2804 0.086905f
C7665 a_42604_n2020 a_46020_n1192 0.043091f
C7666 a_40652_n1572 a_44676_n1572 0.017844f
C7667 a_22052_1944 a_28736_1944 0.019093f
C7668 a_39972_n18440 VDD 0.207295f
C7669 a_23887_n5156 a_24672_n11339 0.020609f
C7670 a_43196_n16916 a_43084_n17349 0.026339f
C7671 a_45660_332 a_42604_n2020 0.064491f
C7672 a_30616_n6221 a_30740_n7464 0.054949f
C7673 a_46916_n18440 a_47004_n18484 0.285629f
C7674 a_45212_n18484 a_45660_n18484 0.012552f
C7675 a_43980_n7941 a_44340_n7844 0.087066f
C7676 a_36724_n7844 a_37172_n7844 0.013276f
C7677 a_41628_n2804 VDD 0.314361f
C7678 a_37484_n9509 a_37844_n9412 0.087174f
C7679 a_23564_n8292 a_24152_n11680 0.028267f
C7680 a_34350_n10980 a_33364_n11384 0.014303f
C7681 a_36588_n11077 a_36500_n10980 0.285629f
C7682 a_43980_n11077 a_44428_n11077 0.012882f
C7683 a_39724_n9509 VDD 0.319134f
C7684 a_28300_n15348 a_27496_n14116 0.028211f
C7685 a_27032_51 VDD 0.244331f
C7686 a_33488_n12996 VDD 0.450166f
C7687 a_21916_n1975 a_27706_n1572 0.023703f
C7688 a_47900_n13780 a_48012_n14213 0.026339f
C7689 a_34796_n14213 a_35244_n14213 0.012882f
C7690 a_33452_n15781 VDD 0.304437f
C7691 a_42076_n2804 a_42188_n3237 0.026339f
C7692 a_24631_n3588 a_22820_n2804 0.145173f
C7693 a_25084_1564 a_22096_376 0.033156f
C7694 a_22500_n1976 a_27736_1248 0.04499f
C7695 a_23932_n18917 VDD 0.302439f
C7696 a_31212_n17349 a_31124_n17252 0.285629f
C7697 a_41740_n17349 a_42188_n17349 0.012882f
C7698 a_47452_n4372 a_47564_n4805 0.026339f
C7699 a_44540_n18484 a_44428_n18917 0.026339f
C7700 a_43980_n6373 a_43892_n6276 0.285629f
C7701 a_25612_n6679 a_29476_n6980 0.086814f
C7702 a_37820_n20052 a_38268_n20052 0.012882f
C7703 a_41764_n20008 a_41852_n20052 0.285629f
C7704 a_43892_n6276 VDD 0.210071f
C7705 a_47116_n11077 a_47028_n10980 0.285629f
C7706 a_28927_n10160 a_31789_n12996 0.075696f
C7707 a_46132_n9412 VDD 0.210512f
C7708 a_41292_n12645 a_41652_n12548 0.087066f
C7709 a_37620_n12548 VDD 0.213356f
C7710 a_37036_n14213 a_37396_n14116 0.087066f
C7711 a_32860_n2020 a_33375_n1976 0.011205f
C7712 a_37844_n15684 VDD 0.214349f
C7713 a_41292_n15781 a_41204_n15684 0.285629f
C7714 a_23564_n20836 a_23844_n16872 0.039686f
C7715 a_45772_n18917 VDD 0.321879f
C7716 a_29332_1243 a_28836_376 0.153696f
C7717 a_42188_n17349 a_42548_n17252 0.087066f
C7718 a_43084_n4805 a_43532_n4805 0.012882f
C7719 a_26956_n18917 a_27316_n18820 0.087066f
C7720 a_22052_n6980 a_22812_n7376 0.011851f
C7721 a_22464_n7393 a_23324_n7420 0.882105f
C7722 a_40172_n18917 a_40620_n18917 0.012001f
C7723 a_47364_n20008 a_47004_n20052 0.086742f
C7724 a_25412_n8501 a_25860_n9032 0.203503f
C7725 a_44340_n3140 VDD 0.212126f
C7726 a_25020_n11383 a_35392_n10172 0.058191f
C7727 a_24965_n9860 a_24684_n16432 0.01818f
C7728 a_23564_n8292 a_21872_n12530 0.021744f
C7729 a_42476_1515 VDD 0.245539f
C7730 a_30871_n11728 VDD 0.96956f
C7731 a_48012_n14213 a_47924_n14116 0.285629f
C7732 a_32308_n1976 a_34953_n1572 0.364092f
C7733 a_39188_n14116 a_39636_n14116 0.013276f
C7734 a_28752_n15348 a_27988_n20388 0.037753f
C7735 a_22500_n1976 a_24128_n704 0.01171f
C7736 a_31684_n16872 VDD 0.215391f
C7737 a_47564_n3237 a_48012_n3237 0.012882f
C7738 a_23564_n17700 a_23484_n16916 0.03f
C7739 a_43532_n3237 a_43444_n3140 0.285629f
C7740 a_24631_n3588 a_25237_n4327 0.085385f
C7741 a_40532_n18820 VDD 0.212561f
C7742 a_25524_1243 a_24913_864 0.035598f
C7743 a_48012_n4805 a_47924_n4708 0.285629f
C7744 a_42548_n17252 a_42996_n17252 0.013276f
C7745 a_21792_n7464 a_22052_n6980 0.088508f
C7746 a_31451_n7508 a_31799_n7508 0.633318f
C7747 a_30781_n452 VDD 0.581638f
C7748 a_37932_n18917 a_37844_n18820 0.285629f
C7749 a_24233_n844 VDD 0.502778f
C7750 a_33564_n20485 a_34012_n20485 0.013103f
C7751 a_33015_n4284 VDD 0.802345f
C7752 a_31460_n10116 a_31872_n10529 0.536965f
C7753 a_32579_769 VDD 0.329304f
C7754 a_46108_n7508 VDD 0.318654f
C7755 a_46916_n10600 VDD 0.205962f
C7756 a_43644_n705 a_43885_n452 0.024891f
C7757 a_26563_n12212 a_27316_n14820 0.57016f
C7758 a_26266_n13736 a_26470_n13736 0.499501f
C7759 a_24233_n13388 a_24128_n13248 0.116059f
C7760 a_40652_n1572 a_45772_n101 0.018297f
C7761 a_44452_n13736 VDD 0.219497f
C7762 a_47900_n1669 a_47812_n1572 0.285629f
C7763 a_45684_n4 VDD 0.213563f
C7764 a_38716_n16916 VDD 0.321613f
C7765 a_23484_n16916 a_23932_n16916 0.012222f
C7766 a_26172_n20052 VDD 0.331989f
C7767 a_37859_377 a_40260_n408 0.146693f
C7768 a_23396_n18440 a_23036_n18484 0.087174f
C7769 a_35156_n18820 a_35604_n18820 0.013276f
C7770 a_42100_n9412 CLK 0.020589f
C7771 a_37372_n9076 a_37820_n9076 0.012882f
C7772 a_41764_n9032 a_41404_n9076 0.087066f
C7773 a_34012_n20485 a_33924_n20388 0.285629f
C7774 a_46108_n4372 VDD 0.318654f
C7775 a_45324_n7941 VDD 0.324845f
C7776 a_37284_n12168 a_37732_n12168 0.013276f
C7777 a_38380_n11077 VDD 0.342539f
C7778 a_31664_n13292 a_32152_n13692 0.08126f
C7779 a_27820_n16432 a_29479_n13735 0.265384f
C7780 a_29161_n14476 VDD 0.484471f
C7781 a_34953_n1572 a_34649_n2412 0.016519f
C7782 a_22820_n2804 a_27452_n2716 0.040289f
C7783 a_42244_n1572 a_42884_n2760 0.038674f
C7784 a_34708_n15304 a_35156_n15304 0.013276f
C7785 a_36140_n17349 VDD 0.313885f
C7786 a_33924_n16872 a_33564_n16916 0.086905f
C7787 a_27988_n20388 a_28076_n18484 0.012909f
C7788 a_22052_n4708 a_22544_n4690 0.015425f
C7789 a_27572_860 a_23004_n2332 0.203342f
C7790 a_39972_n20008 VDD 0.207295f
C7791 a_31236_n18440 a_31684_n18440 0.013276f
C7792 a_43892_n17252 a_44004_n18440 0.026657f
C7793 a_47476_n4708 a_47364_n5896 0.026657f
C7794 a_23887_n5156 a_23324_n7420 0.045083f
C7795 a_25972_n6276 a_31919_n9032 0.037814f
C7796 a_43644_n7508 a_44092_n7508 0.012882f
C7797 a_46916_n9032 a_46556_n9076 0.086742f
C7798 a_44988_n20485 a_45348_n20388 0.087174f
C7799 a_33924_n20388 a_34372_n20388 0.013276f
C7800 a_25831_n11428 a_31565_n9860 0.018657f
C7801 a_41404_n10644 a_41852_n10644 0.012882f
C7802 a_22568_n8944 VDD 0.362583f
C7803 a_44004_n12168 a_43644_n12212 0.087066f
C7804 a_44340_n10980 VDD 0.212126f
C7805 a_46243_769 a_46220_n101 0.029772f
C7806 a_26470_n13736 a_26532_n14437 0.061251f
C7807 a_25132_n16432 a_23608_n15260 1.13433f
C7808 a_39076_n13736 a_39524_n13736 0.013276f
C7809 a_30104_n1148 a_28456_n364 0.061425f
C7810 a_33812_n14116 VDD 0.203482f
C7811 a_31412_n2276 a_31392_n2760 0.573565f
C7812 a_22948_n14820 a_24752_n16132 0.032942f
C7813 a_36948_n17252 VDD 0.21223f
C7814 a_40868_n16872 a_41316_n16872 0.013276f
C7815 a_37284_n16872 a_37372_n16916 0.285629f
C7816 a_43644_n705 a_45660_332 0.01679f
C7817 a_30372_376 a_30104_n1148 0.04944f
C7818 a_26844_n20485 VDD 0.339206f
C7819 a_27988_n4328 a_27485_n10068 0.013149f
C7820 a_41516_n5940 a_41964_n5940 0.013103f
C7821 a_25627_n452 VDD 0.463037f
C7822 a_28324_n20008 a_28772_n20008 0.013276f
C7823 a_22712_n7420 a_25412_n8501 0.022855f
C7824 a_24740_n20008 a_24828_n20052 0.285629f
C7825 a_42748_n10644 CLK 0.012909f
C7826 a_47452_n1669 VDD 0.296789f
C7827 a_41404_n9076 a_41292_n9509 0.026339f
C7828 a_47028_n4708 VDD 0.206217f
C7829 a_30871_n11728 a_32158_n12212 0.033322f
C7830 a_37372_n10644 a_37484_n11077 0.026339f
C7831 a_39972_n9032 VDD 0.207563f
C7832 a_42212_n16872 CLK 0.037136f
C7833 a_47004_n12212 a_47452_n12212 0.012222f
C7834 a_39308_n452 a_39357_n660 0.034588f
C7835 a_27404_n14990 VDD 0.191274f
C7836 a_42300_n15348 a_42748_n15348 0.012882f
C7837 a_24828_n18484 VDD 0.31562f
C7838 a_28144_n4708 a_28548_n5112 0.016877f
C7839 a_43644_n4372 a_44092_n4372 0.012552f
C7840 a_22052_n4708 a_22016_n5825 0.01176f
C7841 a_26756_n20388 VDD 0.204877f
C7842 a_38951_420 a_40776_770 0.34481f
C7843 a_39544_420 a_39352_464 0.934191f
C7844 a_41316_n18440 a_41404_n18484 0.285629f
C7845 a_37372_n18484 a_37820_n18484 0.012882f
C7846 a_39500_n7941 a_39948_n7941 0.012222f
C7847 a_23479_n5156 a_24964_n14116 0.028788f
C7848 a_33497_n9032 a_32767_n9010 0.230761f
C7849 a_42772_n5896 VDD 0.208971f
C7850 a_46556_n10644 a_46668_n11077 0.026339f
C7851 a_22264_n10556 VDD 0.381124f
C7852 a_28232_n12606 a_28040_n12493 0.934191f
C7853 a_44540_n12212 VDD 0.353322f
C7854 a_44452_n15304 VDD 0.219497f
C7855 a_46916_n2760 a_47364_n2760 0.013276f
C7856 a_45572_n2760 a_45660_n2804 0.285629f
C7857 a_21692_n15781 a_22052_n15684 0.086905f
C7858 a_40508_n15348 a_40620_n15781 0.026339f
C7859 a_42604_n2020 a_45572_n1192 0.012511f
C7860 a_40652_n1572 a_44228_n1572 0.016948f
C7861 a_22052_1944 a_22500_n1976 0.019318f
C7862 a_39524_n18440 VDD 0.209499f
C7863 a_23479_n5156 a_24672_n11339 0.038581f
C7864 a_30316_n17349 a_30764_n17349 0.013103f
C7865 a_30616_n6221 a_31068_n6276 0.026665f
C7866 a_46916_n18440 a_46556_n18484 0.086742f
C7867 a_34460_n20052 a_34908_n20052 0.012882f
C7868 a_43980_n7941 a_43892_n7844 0.285629f
C7869 a_25972_n6276 a_28335_n10644 0.048687f
C7870 a_41180_n2804 VDD 0.314361f
C7871 a_44876_n9509 a_45324_n9509 0.012882f
C7872 a_37484_n9509 a_37396_n9412 0.285629f
C7873 a_7119_4292 VDD 1.41434f
C7874 a_39276_n9509 VDD 0.320782f
C7875 a_38604_n12645 a_39052_n12645 0.012552f
C7876 a_31760_n12168 a_33280_n13248 0.097575f
C7877 a_32413_n12996 VDD 0.785627f
C7878 a_38380_n15781 a_38828_n15781 0.012882f
C7879 a_27932_n3543 a_25600_n5895 0.047241f
C7880 a_22820_n2804 a_32359_n4372 0.061452f
C7881 a_25084_1564 a_25936_1564 0.018888f
C7882 a_23484_n18917 VDD 0.301477f
C7883 a_30764_n17349 a_31124_n17252 0.087174f
C7884 a_29196_n18917 a_29644_n18917 0.012882f
C7885 a_43532_n6373 a_43892_n6276 0.087066f
C7886 a_25972_n6276 a_26719_n7464 0.010933f
C7887 a_41764_n20008 a_41404_n20052 0.087066f
C7888 a_47476_n7844 a_47924_n7844 0.013276f
C7889 a_27224_n62 a_28352_n320 0.048436f
C7890 a_29560_n3544 VDD 0.047418f
C7891 a_29992_n11150 a_30808_n10116 0.108733f
C7892 a_32581_n9860 a_31460_n10116 0.025376f
C7893 a_43444_n6276 VDD 0.208665f
C7894 a_46668_n11077 a_47028_n10980 0.087066f
C7895 a_38740_n10980 a_39188_n10980 0.013276f
C7896 a_45684_n9412 VDD 0.212747f
C7897 a_41292_n12645 a_41204_n12548 0.285629f
C7898 a_37172_n12548 VDD 0.211229f
C7899 a_37036_n14213 a_36948_n14116 0.285629f
C7900 a_32636_n2020 a_33375_n1976 0.014035f
C7901 a_45324_n14213 a_45772_n14213 0.012882f
C7902 a_47900_n1236 a_47900_n1669 0.05841f
C7903 a_37396_n15684 VDD 0.211702f
C7904 a_36217_n3500 a_22052_n4708 0.017071f
C7905 a_40620_n15781 a_41204_n15684 0.016748f
C7906 a_29332_1243 a_29744_1564 0.536965f
C7907 a_45324_n18917 VDD 0.324845f
C7908 a_42188_n17349 a_42100_n17252 0.285629f
C7909 a_31124_n17252 a_31572_n17252 0.013276f
C7910 a_38733_n5431 CLK 0.022117f
C7911 a_22464_n7393 a_22712_n7420 0.356609f
C7912 a_26956_n18917 a_26868_n18820 0.285629f
C7913 a_22052_n6980 a_23324_n7420 0.05539f
C7914 a_45212_n20052 a_45660_n20052 0.012552f
C7915 a_41204_n7844 a_41316_n9032 0.026657f
C7916 a_21872_n9394 a_25573_n12167 0.021162f
C7917 a_46916_n20008 a_47004_n20052 0.285629f
C7918 a_43892_n3140 VDD 0.210071f
C7919 a_41864_1394 VDD 1.0704f
C7920 a_23564_n8292 a_23619_n12996 0.042324f
C7921 a_33497_n9032 VDD 0.511582f
C7922 a_22352_n12097 a_22904_n12080 0.361958f
C7923 a_22600_n12124 a_22700_n12080 0.083421f
C7924 VDD VIN 1.54652f
C7925 a_35392_n10172 VDD 0.52824f
C7926 a_42996_n12548 a_43444_n12548 0.013276f
C7927 a_41292_n1669 a_41684_n1976 0.127264f
C7928 a_32736_n1572 a_32100_n1976 0.027448f
C7929 a_47564_n14213 a_47924_n14116 0.087066f
C7930 a_31236_n16872 VDD 0.223727f
C7931 a_42996_n15684 a_43444_n15684 0.013276f
C7932 a_43084_n3237 a_43444_n3140 0.087066f
C7933 a_25237_n4327 a_32359_n4372 0.035939f
C7934 a_35064_1506 a_36192_1248 0.048436f
C7935 a_40084_n18820 VDD 0.207325f
C7936 a_47564_n4805 a_47924_n4708 0.087066f
C7937 a_41652_n4708 a_42100_n4708 0.013276f
C7938 a_23844_n18820 a_24292_n18820 0.013276f
C7939 a_37484_n18917 a_37844_n18820 0.087066f
C7940 a_28352_n320 VDD 0.010384f
C7941 a_47924_n7844 a_47812_n9032 0.026657f
C7942 a_34092_n9076 a_25831_n11428 0.145217f
C7943 a_33120_n3884 VDD 1.78075f
C7944 a_28435_n10599 a_32424_n10512 0.019395f
C7945 a_45660_n7508 VDD 0.320877f
C7946 a_43444_n10980 a_43556_n12168 0.026657f
C7947 a_32854_n12168 a_33686_n11592 0.106585f
C7948 a_40652_n1572 a_45324_n101 0.04743f
C7949 a_46468_n10600 VDD 0.209055f
C7950 a_44004_n13736 VDD 0.2108f
C7951 a_22052_n15304 a_22140_n15348 0.285629f
C7952 a_47452_n1669 a_47812_n1572 0.086635f
C7953 a_42412_n101 a_42324_n4 0.285629f
C7954 a_38268_n16916 VDD 0.356784f
C7955 a_25724_n20052 VDD 0.33355f
C7956 a_22948_n18440 a_23036_n18484 0.285629f
C7957 a_22016_n5825 a_23816_n5408 0.510371f
C7958 a_40420_n7464 a_40868_n7464 0.013276f
C7959 a_33564_n20485 a_33924_n20388 0.087174f
C7960 a_44540_n20485 a_44988_n20485 0.013103f
C7961 a_41316_n9032 a_41404_n9076 0.285629f
C7962 a_43644_n705 EOC 0.01787f
C7963 a_45660_n4372 VDD 0.320877f
C7964 a_38180_n10600 a_38628_n10600 0.013276f
C7965 a_40672_864 VDD 0.010384f
C7966 a_44876_n7941 VDD 0.360805f
C7967 a_37932_n11077 VDD 0.327674f
C7968 a_30903_n13780 a_31455_n13648 0.119687f
C7969 a_31664_n13292 a_31559_n13692 0.536965f
C7970 a_28744_n14432 VDD 1.33211f
C7971 a_23507_n2759 a_25547_n2445 0.010169f
C7972 a_35692_n17349 VDD 0.313885f
C7973 a_27988_n20388 a_27628_n18484 0.051132f
C7974 a_33476_n16872 a_33564_n16916 0.285629f
C7975 a_39524_n20008 VDD 0.209499f
C7976 a_37284_n5896 a_37732_n5896 0.013276f
C7977 a_24492_n5156 a_22464_n7393 0.020315f
C7978 a_23479_n5156 a_23324_n7420 0.02067f
C7979 a_25972_n6276 a_30900_n9032 0.014373f
C7980 a_45684_n18820 a_46132_n18820 0.013276f
C7981 a_25831_n11428 a_29992_n11150 0.046117f
C7982 a_44988_n20485 a_44900_n20388 0.285629f
C7983 a_46468_n9032 a_46556_n9076 0.285629f
C7984 a_31460_n10116 a_31961_n11340 0.043365f
C7985 a_22364_n8944 VDD 0.010384f
C7986 a_39164_n12212 a_39612_n12212 0.012882f
C7987 a_43556_n12168 a_43644_n12212 0.285629f
C7988 a_43892_n10980 VDD 0.210071f
C7989 a_25132_n16432 a_23360_n15233 0.046768f
C7990 a_25831_n12996 a_25160_n14816 0.050403f
C7991 a_33364_n14116 VDD 0.224235f
C7992 a_22948_n14820 a_24088_n16087 0.032681f
C7993 a_27988_n4328 a_22052_n4708 0.051128f
C7994 a_39076_n15304 a_39524_n15304 0.013276f
C7995 a_30555_n2729 a_31392_n2760 0.250931f
C7996 a_31324_n4372 a_32100_n1976 0.104687f
C7997 a_36500_n17252 VDD 0.207483f
C7998 a_40868_n4328 a_41316_n4328 0.013276f
C7999 a_33608_n4284 a_34736_n3840 0.048436f
C8000 a_21604_n3844 a_23887_n5156 0.010754f
C8001 a_29812_860 a_30104_n1148 0.01286f
C8002 a_26396_n20485 VDD 0.330434f
C8003 a_43644_n705 a_45212_332 0.028771f
C8004 a_34012_n18484 a_34460_n18484 0.012882f
C8005 a_24740_n20008 a_24380_n20052 0.087066f
C8006 a_22712_n7420 a_22772_n8944 0.015881f
C8007 a_41852_n7508 a_41740_n7941 0.026339f
C8008 a_26973_n8292 a_27597_n8292 0.104193f
C8009 a_137_4292 a_n199_2852 0.26311f
C8010 a_47004_n1669 VDD 0.296789f
C8011 a_42300_n10644 CLK 0.048577f
C8012 a_44900_n20388 a_45348_n20388 0.013276f
C8013 a_46580_n4708 VDD 0.209016f
C8014 a_24965_n9860 a_23949_n12996 0.021332f
C8015 a_21772_n9860 a_26635_n12996 0.037556f
C8016 a_39524_n9032 VDD 0.209768f
C8017 a_31760_n12168 VDD 0.474597f
C8018 a_41852_n13780 a_42300_n13780 0.012882f
C8019 a_25160_n14816 VDD 1.3448f
C8020 a_37221_n3543 a_39412_n3140 0.015923f
C8021 a_33452_n15348 a_33452_n15781 0.05841f
C8022 a_42884_n2760 a_43332_n2760 0.013276f
C8023 a_24380_n18484 VDD 0.315498f
C8024 a_25600_n5895 a_25412_n5895 0.092015f
C8025 a_43644_n16916 a_44092_n16916 0.012882f
C8026 a_35804_n16916 a_35692_n17349 0.026339f
C8027 a_38951_420 a_39352_464 0.882105f
C8028 a_39056_820 a_40776_770 0.110194f
C8029 a_26308_n20388 VDD 0.205316f
C8030 a_41316_n18440 a_40956_n18484 0.087066f
C8031 a_25972_n6276 a_28624_n9394 0.015298f
C8032 a_31236_n20008 a_31684_n20008 0.013276f
C8033 a_33497_n9032 a_32543_n9032 0.013823f
C8034 a_28454_n2424 VDD 0.690713f
C8035 a_29992_n11150 a_31565_n9860 0.02414f
C8036 a_42324_n5896 VDD 0.208971f
C8037 a_27639_n12537 a_28040_n12493 0.882105f
C8038 a_44540_n12212 a_44428_n12645 0.026339f
C8039 a_44092_n12212 VDD 0.3211f
C8040 a_38268_n13780 a_38380_n14213 0.026339f
C8041 a_45572_n1192 a_46020_n1192 0.013276f
C8042 a_29444_n708 a_31348_n1931 0.026333f
C8043 a_44004_n15304 VDD 0.2108f
C8044 a_45572_n2760 a_45212_n2804 0.086905f
C8045 a_21692_n15781 a_21604_n15684 0.285629f
C8046 a_40652_n1572 a_43780_n1572 0.016172f
C8047 a_39076_n18440 VDD 0.211414f
C8048 a_21692_2431 a_28736_1944 1.14398f
C8049 a_42748_n16916 a_42636_n17349 0.026339f
C8050 a_21792_n7464 a_22264_n5852 0.209412f
C8051 a_45212_332 a_45660_332 0.012222f
C8052 a_46468_n18440 a_46556_n18484 0.285629f
C8053 a_30808_n6334 a_30740_n7464 0.033486f
C8054 a_36276_n7844 a_36724_n7844 0.013276f
C8055 a_43532_n7941 a_43892_n7844 0.087066f
C8056 a_40732_n2804 VDD 0.329307f
C8057 a_26470_n9322 a_26861_n10135 0.032331f
C8058 a_37036_n9509 a_37396_n9412 0.087174f
C8059 a_3025_2852 VDD 1.10914f
C8060 a_34350_n10980 a_28300_n15348 0.091822f
C8061 a_43532_n11077 a_43980_n11077 0.012882f
C8062 a_38828_n9509 VDD 0.323023f
C8063 a_28300_n15348 a_27804_n14165 0.02874f
C8064 a_31789_n12996 VDD 0.594935f
C8065 a_47452_n13780 a_47564_n14213 0.026339f
C8066 a_34348_n14213 a_34796_n14213 0.012882f
C8067 a_28568_n16066 VDD 0.653195f
C8068 a_41628_n2804 a_41740_n3237 0.026339f
C8069 a_23036_n18917 VDD 0.299875f
C8070 a_41292_n17349 a_41740_n17349 0.012882f
C8071 a_30764_n17349 a_30676_n17252 0.285629f
C8072 a_47004_n4372 a_47116_n4805 0.026339f
C8073 a_44092_n18484 a_43980_n18917 0.026339f
C8074 a_43532_n6373 a_43444_n6276 0.285629f
C8075 a_25972_n6276 a_26095_n7464 0.064339f
C8076 a_27032_51 a_27484_n4 0.026665f
C8077 a_37372_n20052 a_37820_n20052 0.012882f
C8078 a_41316_n20008 a_41404_n20052 0.285629f
C8079 a_32189_n9860 a_31460_n10116 0.071389f
C8080 a_40084_n9412 a_40532_n9412 0.013276f
C8081 a_48012_n9509 a_47924_n9412 0.285629f
C8082 a_42412_n101 a_42860_n101 0.012222f
C8083 a_25524_1243 VDD 1.85308f
C8084 a_42996_n6276 VDD 0.205948f
C8085 a_46668_n11077 a_46580_n10980 0.285629f
C8086 a_28927_n10160 a_30340_n12548 0.045344f
C8087 a_40196_1944 OUT[3] 0.021394f
C8088 a_45236_n9412 VDD 0.229781f
C8089 a_36724_n12548 VDD 0.212453f
C8090 a_36588_n14213 a_36948_n14116 0.087066f
C8091 a_32636_n2020 a_32860_n2020 0.066825f
C8092 a_25132_n16432 a_25544_n16412 0.014488f
C8093 a_40652_n1572 OUT[5] 0.010866f
C8094 a_36948_n15684 VDD 0.21223f
C8095 a_40620_n15781 a_40532_n15684 0.285629f
C8096 a_28153_1204 a_28836_376 0.042949f
C8097 a_44876_n18917 VDD 0.360805f
C8098 a_27988_n20388 a_27964_n20052 0.043119f
C8099 a_27988_n4328 a_25573_n12167 0.051242f
C8100 a_41740_n17349 a_42100_n17252 0.087066f
C8101 a_42636_n4805 a_43084_n4805 0.012882f
C8102 a_38403_n5503 CLK 0.018981f
C8103 a_22052_n6980 a_22712_n7420 0.094769f
C8104 a_26508_n18917 a_26868_n18820 0.087066f
C8105 a_39724_n18917 a_40172_n18917 0.012882f
C8106 a_46916_n20008 a_46556_n20052 0.086742f
C8107 a_27485_n8500 a_25573_n12167 0.079847f
C8108 a_43444_n3140 VDD 0.208665f
C8109 a_41616_1564 VDD 0.801558f
C8110 a_36500_n10980 a_36612_n12168 0.026657f
C8111 a_22352_n12097 a_22700_n12080 0.401636f
C8112 a_21940_n11684 a_22904_n12080 0.08126f
C8113 a_33672_n10112 VDD 1.32807f
C8114 a_38740_n14116 a_39188_n14116 0.013276f
C8115 a_32308_n1976 a_32100_n1976 0.426759f
C8116 a_47564_n14213 a_47476_n14116 0.285629f
C8117 a_25647_n1976 a_25547_n2445 0.043074f
C8118 a_22500_n1976 a_27279_n1170 0.022086f
C8119 a_30788_n16872 VDD 0.209936f
C8120 a_25600_n5895 a_28144_n4708 0.101934f
C8121 a_25237_n4327 a_31787_n3969 0.012923f
C8122 a_47116_n3237 a_47564_n3237 0.012882f
C8123 a_43084_n3237 a_42996_n3140 0.285629f
C8124 a_34471_1575 a_36192_1248 0.401636f
C8125 a_39636_n18820 VDD 0.210224f
C8126 a_42100_n17252 a_42548_n17252 0.013276f
C8127 a_47564_n4805 a_47476_n4708 0.285629f
C8128 a_37484_n18917 a_37396_n18820 0.285629f
C8129 a_30451_n452 VDD 0.31647f
C8130 a_29123_n6679 a_31011_n8292 0.035344f
C8131 a_33116_n20485 a_33564_n20485 0.013103f
C8132 a_31460_n10116 a_30808_n10116 0.174595f
C8133 a_24631_n3588 VDD 1.85222f
C8134 a_45212_n7508 VDD 0.342281f
C8135 a_46020_n10600 VDD 0.210736f
C8136 a_40652_n1572 a_42948_n1976 0.025764f
C8137 a_22568_n13648 a_22772_n13648 0.66083f
C8138 a_25642_n13736 a_26266_n13736 0.107109f
C8139 a_43556_n13736 VDD 0.209225f
C8140 a_47452_n1669 a_47364_n1572 0.285629f
C8141 a_22052_n15304 a_21692_n15348 0.086742f
C8142 a_37859_377 a_41533_n727 0.081146f
C8143 a_41336_n407 a_42324_n4 0.010419f
C8144 a_37820_n16916 VDD 0.322978f
C8145 a_23036_n16916 a_23484_n16916 0.012222f
C8146 a_25276_n20052 VDD 0.335085f
C8147 a_22948_n18440 a_22588_n18484 0.087174f
C8148 a_21604_n5412 a_23816_n5408 0.042802f
C8149 a_22364_n5808 a_22568_n5808 0.048436f
C8150 a_22016_n5825 a_24233_n5548 0.020455f
C8151 a_36500_n17252 a_36612_n18440 0.026657f
C8152 a_39524_n4708 a_39357_n5364 0.010897f
C8153 a_27988_n4328 a_27302_n9816 0.014278f
C8154 a_39412_n6276 CLK 0.082282f
C8155 a_34708_n18820 a_35156_n18820 0.013276f
C8156 a_41316_n9032 a_40956_n9076 0.087066f
C8157 a_33564_n20485 a_33476_n20388 0.285629f
C8158 a_27485_n8500 a_27302_n9816 0.017477f
C8159 a_45212_n4372 VDD 0.342281f
C8160 a_44428_n7941 VDD 0.321554f
C8161 a_36700_n12212 a_37284_n12168 0.016748f
C8162 a_35940_2475 OUT[1] 0.023343f
C8163 a_37484_n11077 VDD 0.322148f
C8164 a_27700_n14116 VDD 0.298894f
C8165 a_27316_n14820 a_27524_n15304 0.013419f
C8166 a_22164_n2760 a_23319_n2759 0.101537f
C8167 a_34260_n15304 a_34708_n15304 0.013276f
C8168 a_44340_n14116 a_44452_n15304 0.026657f
C8169 a_23507_n2759 a_24771_n2804 0.015996f
C8170 a_35244_n17349 VDD 0.313885f
C8171 a_22052_n4708 a_22444_n5156 0.122097f
C8172 a_27988_n20388 a_27180_n18484 0.013085f
C8173 a_33476_n16872 a_33116_n16916 0.087174f
C8174 a_39076_n20008 VDD 0.211414f
C8175 a_43444_n17252 a_43556_n18440 0.026657f
C8176 a_30788_n18440 a_31236_n18440 0.013276f
C8177 a_47028_n4708 a_46916_n5896 0.026657f
C8178 a_23887_n5156 a_22464_n7393 0.029087f
C8179 a_43196_n7508 a_43644_n7508 0.012882f
C8180 a_25831_n11428 a_25724_n14564 0.402271f
C8181 a_46468_n9032 a_46108_n9076 0.086905f
C8182 a_33476_n20388 a_33924_n20388 0.013276f
C8183 a_44540_n20485 a_44900_n20388 0.087174f
C8184 a_40956_n10644 a_41404_n10644 0.012882f
C8185 a_31460_n10116 a_31544_n11296 0.034106f
C8186 a_22876_n8988 VDD 0.246128f
C8187 a_28300_n15348 a_34932_n12548 0.01535f
C8188 a_43556_n12168 a_43196_n12212 0.087066f
C8189 a_43444_n10980 VDD 0.208665f
C8190 a_25831_n12996 a_25577_n14956 0.062942f
C8191 a_25524_n708 a_25732_n1192 0.013419f
C8192 a_38628_n13736 a_39076_n13736 0.013276f
C8193 a_30555_n2729 a_31412_n2276 0.033741f
C8194 a_32020_n2276 a_32984_n2672 0.08126f
C8195 a_22140_n15348 a_22140_n15781 0.05841f
C8196 a_36052_n17252 VDD 0.205948f
C8197 a_33015_n4284 a_34736_n3840 0.401636f
C8198 a_21604_n3844 a_23479_n5156 0.029668f
C8199 a_40420_n16872 a_40868_n16872 0.013276f
C8200 a_25948_n20485 VDD 0.333102f
C8201 a_41068_n5940 a_41516_n5940 0.013103f
C8202 a_27876_n20008 a_28324_n20008 0.013276f
C8203 a_24292_n20008 a_24380_n20052 0.285629f
C8204 a_46556_n1669 VDD 0.299954f
C8205 a_41852_n10644 CLK 0.013107f
C8206 a_26470_n9322 a_27302_n9816 0.106585f
C8207 a_46132_n4708 VDD 0.210512f
C8208 a_22264_n8988 a_22016_n13665 0.014653f
C8209 a_21772_n9860 a_26239_n12996 0.09805f
C8210 a_24965_n9860 a_22264_n13692 0.049344f
C8211 a_39076_n9032 VDD 0.211682f
C8212 a_46556_n12212 a_47004_n12212 0.012222f
C8213 a_25577_n14956 VDD 0.481263f
C8214 a_41852_n15348 a_42300_n15348 0.012882f
C8215 a_38996_n408 a_39556_n4 0.302602f
C8216 a_23932_n18484 VDD 0.302439f
C8217 a_43196_n4372 a_43644_n4372 0.012552f
C8218 a_25860_n20388 VDD 0.20723f
C8219 a_39056_820 a_39352_464 0.05539f
C8220 a_40868_n18440 a_40956_n18484 0.285629f
C8221 a_23887_n5156 a_26973_n8292 0.015899f
C8222 a_24672_n11339 a_24752_n8292 0.043704f
C8223 a_23479_n5156 a_27597_n8292 0.023525f
C8224 a_39052_n7941 a_39500_n7941 0.013103f
C8225 a_27452_n2716 VDD 0.281291f
C8226 a_41876_n5896 VDD 0.208971f
C8227 a_46108_n10644 a_46220_n11077 0.026339f
C8228 a_30296_n10980 a_30500_n10980 0.66083f
C8229 a_29744_n10980 a_31856_n11296 0.277491f
C8230 a_45684_n4 a_46132_n4 0.013276f
C8231 a_23619_n9860 VDD 0.318017f
C8232 a_27639_n12537 a_27535_n12493 0.277491f
C8233 a_43644_n12212 VDD 0.319164f
C8234 a_29444_n708 a_27988_n4328 0.030019f
C8235 a_26239_n12996 a_27085_n16132 0.017088f
C8236 a_25132_n16432 a_24752_n16132 0.011963f
C8237 a_43556_n15304 VDD 0.209225f
C8238 a_40060_n15348 a_40172_n15781 0.026339f
C8239 a_46468_n2760 a_46916_n2760 0.013276f
C8240 a_45124_n2760 a_45212_n2804 0.285629f
C8241 a_40652_n1572 a_43332_n1572 0.017033f
C8242 a_21692_2431 a_22500_n1976 0.01978f
C8243 a_38628_n18440 VDD 0.214363f
C8244 a_29868_n17349 a_30316_n17349 0.013103f
C8245 a_22544_n4690 a_24672_n11339 0.029473f
C8246 a_21792_n7464 a_22016_n5825 0.042591f
C8247 a_23479_n5156 a_24492_n5156 1.49671f
C8248 a_30808_n6334 a_31068_n6276 0.66083f
C8249 a_46468_n18440 a_46108_n18484 0.086905f
C8250 a_30215_n6265 a_30740_n7464 0.375982f
C8251 a_43532_n7941 a_43444_n7844 0.285629f
C8252 a_34012_n20052 a_34460_n20052 0.012882f
C8253 a_26266_n9240 a_26861_n10135 0.014311f
C8254 a_44428_n9509 a_44876_n9509 0.012882f
C8255 a_37036_n9509 a_36948_n9412 0.285629f
C8256 a_35064_n11383 a_28300_n15348 0.194175f
C8257 a_34350_n10980 a_34538_n10980 0.025208f
C8258 a_38380_n9509 VDD 0.34331f
C8259 a_38156_n12645 a_38604_n12645 0.012552f
C8260 a_29360_n12864 VDD 0.010384f
C8261 a_27709_n16132 VDD 0.710574f
C8262 a_27932_n3543 a_27337_n3140 0.100784f
C8263 a_37932_n15781 a_38380_n15781 0.012882f
C8264 a_26607_n3544 a_25600_n5895 0.018734f
C8265 a_22588_n18917 VDD 0.296789f
C8266 a_30316_n17349 a_30676_n17252 0.087174f
C8267 a_28748_n18917 a_29196_n18917 0.012882f
C8268 a_22220_n9860 a_22568_n8944 0.017396f
C8269 a_43084_n6373 a_43444_n6276 0.087066f
C8270 a_25972_n6276 a_25685_n7463 0.163589f
C8271 a_24672_n11339 a_21872_n9394 0.027505f
C8272 a_47028_n7844 a_47476_n7844 0.013276f
C8273 a_41316_n20008 a_40956_n20052 0.087066f
C8274 a_31565_n9860 a_31460_n10116 0.02673f
C8275 a_47564_n9509 a_47924_n9412 0.087066f
C8276 a_24628_1252 VDD 0.533626f
C8277 a_42548_n6276 VDD 0.205948f
C8278 a_31544_n11296 a_32026_n12168 0.023072f
C8279 a_46220_n11077 a_46580_n10980 0.087066f
C8280 a_38292_n10980 a_38740_n10980 0.013276f
C8281 a_28927_n10160 a_31459_n12996 0.027135f
C8282 a_44788_n9412 VDD 0.22479f
C8283 a_40396_n12645 a_40308_n12548 0.285629f
C8284 a_36276_n12548 VDD 0.209521f
C8285 a_36588_n14213 a_36500_n14116 0.285629f
C8286 a_44876_n14213 a_45324_n14213 0.012882f
C8287 a_47452_n1236 a_47452_n1669 0.05841f
C8288 a_36500_n15684 VDD 0.207483f
C8289 a_40172_n15781 a_40532_n15684 0.086635f
C8290 a_22948_n15684 a_22948_n16872 0.05841f
C8291 a_44428_n18917 VDD 0.321554f
C8292 a_27988_n20388 a_27516_n20052 0.030501f
C8293 a_41740_n17349 a_41652_n17252 0.285629f
C8294 a_30676_n17252 a_31124_n17252 0.013276f
C8295 a_23479_n5156 a_22568_n5808 0.027985f
C8296 a_22052_n6980 a_22464_n7393 0.536965f
C8297 a_26508_n18917 a_26420_n18820 0.285629f
C8298 a_46468_n20008 a_46556_n20052 0.285629f
C8299 a_42996_n3140 VDD 0.205948f
C8300 a_22352_n12097 a_23212_n12124 0.882105f
C8301 a_21940_n11684 a_22700_n12080 0.011851f
C8302 a_34089_n10252 VDD 0.475141f
C8303 a_42548_n12548 a_42996_n12548 0.013276f
C8304 a_31324_n4372 a_31405_n452 0.054409f
C8305 a_47116_n14213 a_47476_n14116 0.087066f
C8306 a_32308_n1572 a_32100_n1976 0.015646f
C8307 a_22500_n1976 a_27055_n1192 0.012805f
C8308 a_30340_n16872 VDD 0.132142f
C8309 a_27337_n3140 a_27540_n3797 0.03884f
C8310 a_42636_n3237 a_42996_n3140 0.087066f
C8311 a_42548_n15684 a_42996_n15684 0.013276f
C8312 a_39188_n18820 VDD 0.211952f
C8313 a_47116_n4805 a_47476_n4708 0.087066f
C8314 a_41204_n4708 a_41652_n4708 0.013276f
C8315 a_23564_n20836 a_24292_n20008 0.019525f
C8316 a_37036_n18917 a_37396_n18820 0.087066f
C8317 a_44340_n6276 a_44452_n7464 0.026657f
C8318 a_23396_n18820 a_23844_n18820 0.013276f
C8319 a_22220_n9860 a_22264_n10556 0.023052f
C8320 a_28456_n364 VDD 0.384715f
C8321 a_22568_n1104 VDD 0.360568f
C8322 a_47476_n7844 a_47364_n9032 0.026657f
C8323 a_33832_n8572 a_34092_n9076 0.551506f
C8324 a_32359_n4372 VDD 1.30891f
C8325 a_44340_n9412 a_44452_n10600 0.026657f
C8326 a_28435_n10599 a_32732_n10556 0.013768f
C8327 a_30136_n10600 a_30808_n10116 0.037845f
C8328 a_30372_376 VDD 0.605104f
C8329 a_47812_n7464 VDD 0.211703f
C8330 a_42996_n10980 a_43108_n12168 0.026657f
C8331 a_32650_n12168 a_32854_n12168 0.499501f
C8332 a_45572_n10600 VDD 0.213324f
C8333 a_25237_n13735 a_26266_n13736 0.055203f
C8334 a_40652_n1572 a_44509_n452 0.013465f
C8335 a_43108_n13736 VDD 0.206217f
C8336 a_36500_n14116 a_36500_n15304 0.05841f
C8337 a_47004_n1669 a_47364_n1572 0.086742f
C8338 a_21604_n15304 a_21692_n15348 0.285629f
C8339 a_37859_377 a_41203_n799 0.042383f
C8340 a_37372_n16916 VDD 0.324575f
C8341 a_40652_n1572 a_45012_1564 0.01621f
C8342 a_31961_1204 a_32909_841 0.016355f
C8343 a_24828_n20052 VDD 0.349007f
C8344 a_22500_n18440 a_22588_n18484 0.285629f
C8345 a_22876_n5852 a_22568_n5808 0.934191f
C8346 a_25636_n18440 a_26084_n18440 0.013276f
C8347 a_21604_n5412 a_24233_n5548 0.019043f
C8348 a_39972_n7464 a_40420_n7464 0.013276f
C8349 a_48012_n18917 a_47924_n18820 0.285629f
C8350 a_33116_n20485 a_33476_n20388 0.087174f
C8351 a_40868_n9032 a_40956_n9076 0.285629f
C8352 a_47812_n4328 VDD 0.211703f
C8353 a_37732_n10600 a_38180_n10600 0.013276f
C8354 a_43980_n7941 VDD 0.31896f
C8355 a_37036_n11077 VDD 0.334604f
C8356 a_30903_n13780 a_31559_n13692 0.510371f
C8357 a_27496_n14116 VDD 0.360568f
C8358 a_27852_n14990 a_28212_n15303 0.015869f
C8359 a_22164_n2760 a_22672_n2759 0.014431f
C8360 a_41684_n1976 a_41988_n2760 0.018735f
C8361 a_34796_n17349 VDD 0.313885f
C8362 a_22052_n4708 a_21604_n5067 0.197884f
C8363 a_33028_n16872 a_33116_n16916 0.285629f
C8364 a_36164_n16872 a_36612_n16872 0.013276f
C8365 a_38628_n20008 VDD 0.214363f
C8366 a_22444_n5156 a_23016_n7376 0.016397f
C8367 a_23479_n5156 a_22464_n7393 0.039108f
C8368 a_29612_n8292 a_37284_n5896 0.018575f
C8369 a_25972_n6276 a_28617_n8548 0.131328f
C8370 a_45236_n18820 a_45684_n18820 0.013276f
C8371 a_28671_n1976 VDD 0.729619f
C8372 a_44540_n20485 a_44452_n20388 0.285629f
C8373 a_46020_n9032 a_46108_n9076 0.285629f
C8374 a_47364_n9032 a_47812_n9032 0.013276f
C8375 a_42948_n1976 a_43556_n661 0.014295f
C8376 a_22264_n8988 VDD 0.644454f
C8377 a_38716_n12212 a_39164_n12212 0.012882f
C8378 a_24964_n14116 a_27820_n16432 0.104133f
C8379 a_43108_n12168 a_43196_n12212 0.285629f
C8380 a_28300_n15348 a_34484_n12548 0.034232f
C8381 a_42996_n10980 VDD 0.205948f
C8382 a_28736_1944 a_26631_7 0.051948f
C8383 a_38628_n15304 a_39076_n15304 0.013276f
C8384 a_32020_n2276 a_32780_n2672 0.011851f
C8385 a_35604_n17252 VDD 0.205948f
C8386 a_40420_n4328 a_40868_n4328 0.013276f
C8387 a_33120_n3884 a_34736_n3840 0.011851f
C8388 a_43644_n705 a_47197_908 0.466489f
C8389 a_40652_n1572 a_42604_n2020 0.763658f
C8390 a_25500_n20485 VDD 0.341359f
C8391 a_33564_n18484 a_34012_n18484 0.012882f
C8392 a_41404_n7508 a_41292_n7941 0.026339f
C8393 a_24292_n20008 a_23932_n20052 0.087066f
C8394 a_46580_n4 VDD 0.209833f
C8395 a_46108_n1669 VDD 0.300761f
C8396 a_40508_n9076 a_40620_n9509 0.026339f
C8397 a_44452_n20388 a_44900_n20388 0.013276f
C8398 a_45684_n4708 VDD 0.212747f
C8399 a_21772_n9860 a_25831_n12996 0.035249f
C8400 a_22264_n8988 a_21604_n13252 0.013592f
C8401 a_38628_n9032 VDD 0.214632f
C8402 a_30787_n12167 VDD 0.479437f
C8403 a_41404_n13780 a_41852_n13780 0.012882f
C8404 a_38733_n2295 a_37452_n3888 0.0189f
C8405 a_42436_n2760 a_42884_n2760 0.013276f
C8406 a_22820_n2804 a_28583_n3140 0.022917f
C8407 a_39308_n452 a_39556_n4 0.026144f
C8408 a_23484_n18484 VDD 0.301477f
C8409 a_43196_n16916 a_43644_n16916 0.012882f
C8410 a_35356_n16916 a_35244_n17349 0.026339f
C8411 a_25412_n20388 VDD 0.231301f
C8412 a_38951_420 a_38847_464 0.277491f
C8413 a_23479_n5156 a_26973_n8292 0.082782f
C8414 a_40868_n18440 a_40508_n18484 0.087066f
C8415 a_30788_n20008 a_31236_n20008 0.013276f
C8416 a_25895_n2624 VDD 0.240607f
C8417 a_41428_n5896 VDD 0.208971f
C8418 a_30604_n11029 a_31544_n11296 0.056721f
C8419 a_29744_n10980 a_31961_n11340 0.020455f
C8420 a_21772_n9860 VDD 1.04197f
C8421 a_27639_n12537 a_28232_n12606 0.361958f
C8422 a_44092_n12212 a_43980_n12645 0.026339f
C8423 a_43196_n12212 VDD 0.316157f
C8424 a_37820_n13780 a_37932_n14213 0.026339f
C8425 a_45124_n1192 a_45572_n1192 0.013276f
C8426 a_43108_n15304 VDD 0.206217f
C8427 a_22588_n15781 a_23036_n15781 0.012552f
C8428 a_38180_n18440 VDD 0.245127f
C8429 a_23479_n5156 a_23887_n5156 0.042199f
C8430 a_42300_n16916 a_42188_n17349 0.026339f
C8431 a_21792_n7464 a_21604_n5412 0.013914f
C8432 a_46573_841 a_42604_n2020 0.021188f
C8433 a_36700_n18484 a_36588_n18917 0.026339f
C8434 a_30808_n6334 a_30616_n6221 0.934191f
C8435 a_47364_n18440 a_47812_n18440 0.013276f
C8436 a_46020_n18440 a_46108_n18484 0.285629f
C8437 a_43084_n7941 a_43444_n7844 0.087066f
C8438 a_36588_n9509 a_36948_n9412 0.087174f
C8439 a_26266_n9240 a_26531_n10207 0.010173f
C8440 a_137_4292 VIN 0.226767f
C8441 a_25524_n6635 VDD 0.557737f
C8442 a_43084_n11077 a_43532_n11077 0.012882f
C8443 a_23564_n11428 a_22352_n12097 0.028233f
C8444 a_37932_n9509 VDD 0.328094f
C8445 a_28300_n15348 a_26944_n14116 0.02091f
C8446 a_30340_n12548 VDD 0.131135f
C8447 a_33900_n14213 a_34348_n14213 0.012882f
C8448 a_47004_n13780 a_47116_n14213 0.026339f
C8449 a_27085_n16132 VDD 0.586003f
C8450 a_41180_n2804 a_41292_n3237 0.026339f
C8451 a_26383_n2968 a_25600_n5895 0.01183f
C8452 a_23004_n2332 a_22164_n2760 0.109383f
C8453 a_22052_1944 a_28836_376 0.02931f
C8454 a_25084_1564 a_25524_1243 0.026957f
C8455 a_22140_n18917 VDD 0.296789f
C8456 a_30316_n17349 a_30228_n17252 0.285629f
C8457 a_46556_n4372 a_46668_n4805 0.026339f
C8458 a_43644_n18484 a_43532_n18917 0.026339f
C8459 a_43084_n6373 a_42996_n6276 0.285629f
C8460 a_40868_n20008 a_40956_n20052 0.285629f
C8461 a_39636_n9412 a_40084_n9412 0.013276f
C8462 a_47564_n9509 a_47476_n9412 0.285629f
C8463 a_42100_n6276 VDD 0.205948f
C8464 a_46220_n11077 a_46132_n10980 0.285629f
C8465 a_25724_n14564 a_25642_n13736 0.019194f
C8466 a_28927_n10160 a_30428_n12645 0.030982f
C8467 a_44340_n9412 VDD 0.212126f
C8468 a_24684_n16432 a_25160_n14816 0.010208f
C8469 a_39948_n12645 a_40308_n12548 0.086635f
C8470 a_35828_n12548 VDD 0.209521f
C8471 a_36140_n14213 a_36500_n14116 0.087066f
C8472 a_36052_n15684 VDD 0.205948f
C8473 a_40172_n15781 a_40084_n15684 0.285629f
C8474 a_43980_n18917 VDD 0.31896f
C8475 a_42188_n4805 a_42636_n4805 0.012882f
C8476 a_41292_n17349 a_41652_n17252 0.087066f
C8477 a_26060_n18917 a_26420_n18820 0.087066f
C8478 a_39276_n18917 a_39724_n18917 0.012882f
C8479 a_21872_n9394 a_25860_n9032 0.058751f
C8480 a_40308_n7844 a_40420_n9032 0.026657f
C8481 a_46468_n20008 a_46108_n20052 0.086905f
C8482 a_42548_n3140 VDD 0.205948f
C8483 a_22876_n10556 a_23816_n10112 0.056721f
C8484 a_32856_n7376 VDD 0.244843f
C8485 a_22352_n12097 a_22600_n12124 0.355778f
C8486 a_32158_n12212 a_30787_n12167 0.012593f
C8487 a_21940_n11684 a_23212_n12124 0.05539f
C8488 a_47116_n14213 a_47028_n14116 0.285629f
C8489 a_38292_n14116 a_38740_n14116 0.013276f
C8490 a_22500_n1976 a_26431_n1192 0.012702f
C8491 a_28636_n16916 VDD 0.327167f
C8492 a_27337_n3140 a_28144_n4708 0.194255f
C8493 a_42636_n3237 a_42548_n3140 0.285629f
C8494 a_46668_n3237 a_47116_n3237 0.012882f
C8495 a_38740_n18820 VDD 0.214614f
C8496 a_23564_n20836 a_23844_n20008 0.038226f
C8497 a_28436_n17252 a_28436_n18440 0.05841f
C8498 a_47116_n4805 a_47028_n4708 0.285629f
C8499 a_41652_n17252 a_42100_n17252 0.013276f
C8500 a_37036_n18917 a_36948_n18820 0.285629f
C8501 a_29123_n6679 a_28764_n8247 0.627026f
C8502 a_22364_n1104 VDD 0.010384f
C8503 a_31787_n3969 VDD 0.673512f
C8504 a_29812_860 VDD 0.540215f
C8505 a_29992_n11150 a_30092_n10980 0.094174f
C8506 a_28435_n10599 a_31872_n10529 0.020772f
C8507 a_47364_n7464 VDD 0.205948f
C8508 a_45124_n10600 VDD 0.26277f
C8509 a_25237_n13735 a_25642_n13736 0.590436f
C8510 a_22876_n13692 a_22772_n13648 0.026665f
C8511 a_42660_n13736 VDD 0.206217f
C8512 a_47004_n1669 a_46916_n1572 0.285629f
C8513 a_44452_n16872 VDD 0.219497f
C8514 a_22588_n16916 a_23036_n16916 0.012552f
C8515 a_40652_n1572 a_43644_n705 0.136576f
C8516 a_24380_n20052 VDD 0.347672f
C8517 a_45100_1467 a_45012_1564 0.285629f
C8518 a_27988_n20388 a_28300_n20485 0.016742f
C8519 a_36052_n17252 a_36164_n18440 0.026657f
C8520 a_22500_n18440 a_22140_n18484 0.087174f
C8521 a_22264_n5852 a_22568_n5808 0.011343f
C8522 a_47564_n18917 a_47924_n18820 0.087066f
C8523 a_34260_n18820 a_34708_n18820 0.013276f
C8524 a_44228_n1192 VDD 0.138446f
C8525 a_33116_n20485 a_33028_n20388 0.285629f
C8526 a_23564_n8292 a_23816_n10112 0.021155f
C8527 a_40868_n9032 a_40508_n9076 0.087066f
C8528 a_47364_n4328 VDD 0.205948f
C8529 a_32581_n9860 a_33364_n11384 0.575258f
C8530 a_25020_n11383 a_34350_n10980 0.403659f
C8531 a_44452_376 VDD 0.138628f
C8532 a_43532_n7941 VDD 0.317216f
C8533 a_36252_n12212 a_36700_n12212 0.012552f
C8534 a_36588_n11077 VDD 0.334684f
C8535 a_30903_n13780 a_31664_n13292 0.042802f
C8536 a_27292_n14116 VDD 0.010384f
C8537 a_34248_n3310 a_33292_n2716 0.010362f
C8538 a_43892_n14116 a_44004_n15304 0.026657f
C8539 a_27404_n14990 a_28212_n15303 0.089794f
C8540 a_24403_n2414 a_24771_n2804 0.514036f
C8541 a_33812_n15304 a_34260_n15304 0.013276f
C8542 a_35849_n1192 a_33077_n1191 0.014677f
C8543 a_34348_n17349 VDD 0.313885f
C8544 a_33028_n16872 a_32668_n16916 0.087174f
C8545 a_23564_n17700 a_28524_n17349 0.030152f
C8546 a_37844_1564 a_38295_332 0.018588f
C8547 a_28492_332 a_28132_376 0.574924f
C8548 a_38180_n20008 VDD 0.245127f
C8549 VDD OUT[1] 1.1452f
C8550 a_46580_n4708 a_46468_n5896 0.026657f
C8551 a_42996_n17252 a_43108_n18440 0.026657f
C8552 a_30340_n18440 a_30788_n18440 0.013276f
C8553 a_42748_n7508 a_43196_n7508 0.012882f
C8554 a_26495_n1976 VDD 0.319963f
C8555 a_33028_n20388 a_33476_n20388 0.013276f
C8556 a_46020_n9032 a_45660_n9076 0.086905f
C8557 a_43868_n20485 a_44452_n20388 0.016748f
C8558 a_40508_n10644 a_40956_n10644 0.012882f
C8559 a_44452_n10600 a_44540_n10644 0.285629f
C8560 a_42948_n1976 a_42972_n1236 0.048279f
C8561 a_22016_n8961 VDD 0.799451f
C8562 a_27281_n16854 a_27852_n14990 0.055894f
C8563 a_43108_n12168 a_42748_n12212 0.087066f
C8564 a_42548_n10980 VDD 0.205948f
C8565 a_38180_n13736 a_38628_n13736 0.013276f
C8566 a_25132_n16432 a_22948_n14820 0.013508f
C8567 a_22500_n1976 a_26631_7 0.04046f
C8568 a_32020_n2276 a_33292_n2716 0.05539f
C8569 a_21692_n15348 a_21692_n15781 0.05841f
C8570 a_35156_n17252 VDD 0.205948f
C8571 a_39972_n16872 a_40420_n16872 0.013276f
C8572 a_21792_n7464 a_22444_n5156 0.064161f
C8573 a_40652_n1572 a_45660_332 0.023143f
C8574 a_43644_n705 a_46573_841 0.089517f
C8575 a_24604_n20485 VDD 0.396125f
C8576 a_40620_n5940 a_41068_n5940 0.013103f
C8577 a_44116_n5896 a_44204_n5940 0.285629f
C8578 a_26643_n8292 a_26973_n8292 0.538085f
C8579 a_22712_n7420 a_21872_n9394 1.08125f
C8580 a_137_4292 a_3025_2852 0.278387f
C8581 a_23844_n20008 a_23932_n20052 0.285629f
C8582 a_27428_n20008 a_27876_n20008 0.013276f
C8583 a_45660_n1669 VDD 0.302997f
C8584 a_45236_n4708 VDD 0.229781f
C8585 a_24965_n9860 a_21872_n12530 0.027365f
C8586 a_38180_n9032 VDD 0.24541f
C8587 a_46108_n12212 a_46556_n12212 0.012552f
C8588 a_47812_n12168 a_47900_n12212 0.285629f
C8589 a_31664_n13292 a_33452_n14213 0.059049f
C8590 a_21604_n708 a_23542_n1754 0.061254f
C8591 a_22164_n2760 a_25600_n5895 0.207267f
C8592 a_38403_n2367 a_37452_n3888 0.215002f
C8593 a_41404_n15348 a_41852_n15348 0.012882f
C8594 a_23004_n2332 a_22918_n2020 0.09006f
C8595 a_39308_n452 a_38996_n408 0.092494f
C8596 a_23036_n18484 VDD 0.299875f
C8597 a_39056_820 a_39556_n4 0.065185f
C8598 a_42748_n4372 a_43196_n4372 0.012552f
C8599 a_38951_420 a_39544_420 0.361958f
C8600 a_38295_332 a_39352_464 0.056721f
C8601 a_24516_n20388 VDD 0.236934f
C8602 a_22444_n5156 a_28764_n8247 0.010541f
C8603 a_23887_n5156 a_26643_n8292 0.214077f
C8604 a_40420_n18440 a_40508_n18484 0.285629f
C8605 a_44004_n18440 a_44452_n18440 0.013276f
C8606 a_38604_n7941 a_39052_n7941 0.013103f
C8607 a_26499_n2732 VDD 0.271393f
C8608 a_40980_n5896 VDD 0.20894f
C8609 a_30604_n11029 a_30500_n10980 0.026665f
C8610 a_30092_n10980 a_30296_n10980 0.048436f
C8611 a_29744_n10980 a_31544_n11296 0.510371f
C8612 a_45660_n10644 a_45772_n11077 0.026339f
C8613 a_34986_n9032 VDD 0.014149f
C8614 a_42748_n12212 VDD 0.315469f
C8615 a_29444_n708 a_30584_n1954 0.065269f
C8616 a_42660_n15304 VDD 0.206217f
C8617 a_46020_n2760 a_46468_n2760 0.013276f
C8618 a_39612_n15348 a_39724_n15781 0.026339f
C8619 a_42604_n2020 a_43556_n661 0.012116f
C8620 a_37732_n18440 VDD 0.213126f
C8621 a_26383_1944 a_26607_1966 0.538085f
C8622 a_35849_n1192 a_35568_n4 0.042968f
C8623 a_29420_n17349 a_29868_n17349 0.013103f
C8624 a_22544_n4690 a_24492_n5156 0.025357f
C8625 a_22444_n5156 a_24672_n11339 0.017941f
C8626 a_46243_769 a_42604_n2020 0.217243f
C8627 a_30215_n6265 a_30616_n6221 0.882105f
C8628 a_46020_n18440 a_45660_n18484 0.086905f
C8629 a_33564_n20052 a_34012_n20052 0.012882f
C8630 a_43084_n7941 a_42996_n7844 0.285629f
C8631 a_43980_n9509 a_44428_n9509 0.012882f
C8632 a_36588_n9509 a_36500_n9412 0.285629f
C8633 a_25612_n6679 VDD 0.661995f
C8634 a_37484_n9509 VDD 0.322568f
C8635 a_37708_n12645 a_38156_n12645 0.012552f
C8636 a_31459_n12996 VDD 0.358583f
C8637 a_21916_n1975 a_26495_n1976 0.021179f
C8638 a_23564_n20836 VDD 1.45885f
C8639 a_37484_n15781 a_37932_n15781 0.012882f
C8640 a_26607_n3544 a_27337_n3140 0.237391f
C8641 a_31324_n4372 a_29560_n3544 0.016211f
C8642 a_21692_n18917 VDD 0.300735f
C8643 a_25084_1564 a_24628_1252 0.308631f
C8644 a_29868_n17349 a_30228_n17252 0.087174f
C8645 a_28300_n18917 a_28748_n18917 0.012882f
C8646 a_22220_n9860 a_22876_n8988 0.017563f
C8647 a_42636_n6373 a_42996_n6276 0.087066f
C8648 a_40868_n20008 a_40508_n20052 0.087066f
C8649 a_46580_n7844 a_47028_n7844 0.013276f
C8650 a_47116_n9509 a_47476_n9412 0.087066f
C8651 a_32581_n9860 a_28435_n10599 0.546444f
C8652 a_41652_n6276 VDD 0.205948f
C8653 a_37844_n10980 a_38292_n10980 0.013276f
C8654 a_25724_n14564 a_25237_n13735 0.302409f
C8655 a_45772_n11077 a_46132_n10980 0.087066f
C8656 a_43892_n9412 VDD 0.210071f
C8657 a_39948_n12645 a_39860_n12548 0.285629f
C8658 a_25132_n16432 a_25642_n13736 0.046405f
C8659 a_24684_n16432 a_25577_n14956 0.013666f
C8660 a_35380_n12548 VDD 0.209521f
C8661 a_36140_n14213 a_36052_n14116 0.285629f
C8662 a_44428_n14213 a_44876_n14213 0.012882f
C8663 a_47004_n1236 a_47004_n1669 0.05841f
C8664 a_35604_n15684 VDD 0.205948f
C8665 a_22500_n15684 a_22500_n16872 0.05841f
C8666 a_39724_n15781 a_40084_n15684 0.087066f
C8667 a_43532_n18917 VDD 0.317216f
C8668 a_41292_n17349 a_41204_n17252 0.285629f
C8669 a_22544_n4690 a_22568_n5808 0.046848f
C8670 a_23479_n5156 a_22876_n5852 0.041865f
C8671 a_23887_n5156 a_22264_n5852 0.010666f
C8672 a_30228_n17252 a_30676_n17252 0.013276f
C8673 a_26060_n18917 a_25972_n18820 0.285629f
C8674 a_47364_n20008 a_47812_n20008 0.013276f
C8675 a_21872_n9394 a_25412_n8501 0.010484f
C8676 a_46020_n20008 a_46108_n20052 0.285629f
C8677 a_42100_n3140 VDD 0.205948f
C8678 a_22016_n10529 a_23816_n10112 0.510371f
C8679 a_21940_n11684 a_22600_n12124 0.098559f
C8680 a_42100_n12548 a_42548_n12548 0.013276f
C8681 a_46668_n14213 a_47028_n14116 0.087066f
C8682 a_37221_n3543 a_40196_n1884 0.565269f
C8683 a_24578_n2020 a_24771_n2804 0.027818f
C8684 a_23564_n17700 a_28548_n16872 0.037833f
C8685 a_42100_n15684 a_42548_n15684 0.013276f
C8686 a_42188_n3237 a_42548_n3140 0.087066f
C8687 a_22096_376 a_22116_860 0.577309f
C8688 a_34576_1204 a_36192_1248 0.011851f
C8689 a_38292_n18820 VDD 0.244791f
C8690 a_46668_n4805 a_47028_n4708 0.087066f
C8691 a_22948_n18820 a_23396_n18820 0.013276f
C8692 a_36588_n18917 a_36948_n18820 0.087066f
C8693 a_43892_n6276 a_44004_n7464 0.026657f
C8694 a_22876_n1148 VDD 0.243199f
C8695 a_47028_n7844 a_46916_n9032 0.026657f
C8696 a_43892_n9412 a_44004_n10600 0.026657f
C8697 a_46916_n7464 VDD 0.205962f
C8698 a_32026_n12168 a_32650_n12168 0.107109f
C8699 a_42548_n10980 a_42660_n12168 0.026657f
C8700 a_44540_n10644 VDD 0.353322f
C8701 a_26239_n12996 a_27192_n14286 0.016811f
C8702 a_42212_n13736 VDD 0.206217f
C8703 a_21604_n15304 a_22052_n15304 0.013276f
C8704 a_27988_n4328 a_31392_n2760 0.051379f
C8705 a_36052_n14116 a_36052_n15304 0.05841f
C8706 a_46556_n1669 a_46916_n1572 0.086742f
C8707 a_44004_n16872 VDD 0.2108f
C8708 a_45100_1467 a_43644_n705 0.015159f
C8709 a_37859_377 a_39352_464 0.043558f
C8710 a_23932_n20052 VDD 0.318353f
C8711 a_25188_n18440 a_25636_n18440 0.013276f
C8712 a_27988_n20388 a_27540_n20747 0.225775f
C8713 a_22444_n5156 a_30740_n7464 0.014258f
C8714 a_22052_n18440 a_22140_n18484 0.285629f
C8715 a_22264_n5852 a_22364_n5808 0.094469f
C8716 a_38628_n4708 a_38733_n5431 0.040915f
C8717 a_22016_n5825 a_22568_n5808 0.361958f
C8718 a_22712_n7420 a_23564_n8292 0.03498f
C8719 a_39524_n7464 a_39972_n7464 0.013276f
C8720 a_47564_n18917 a_47476_n18820 0.285629f
C8721 a_42884_n1192 VDD 0.125706f
C8722 a_43420_n20485 a_43868_n20485 0.013103f
C8723 a_40420_n9032 a_40508_n9076 0.285629f
C8724 a_32444_n20485 a_33028_n20388 0.016748f
C8725 a_46916_n4328 VDD 0.205962f
C8726 a_40260_n408 VDD 0.67476f
C8727 a_37284_n10600 a_37732_n10600 0.013276f
C8728 a_25020_n11383 a_35064_n11383 0.052712f
C8729 a_43084_n7941 VDD 0.313885f
C8730 a_34350_n10980 VDD 0.366554f
C8731 a_30159_n13296 a_29479_n13735 0.184288f
C8732 a_27804_n14165 VDD 0.243827f
C8733 a_22820_n2804 a_22672_n2759 0.150657f
C8734 a_33900_n17349 VDD 0.313885f
C8735 a_35716_n16872 a_36164_n16872 0.013276f
C8736 a_32580_n16872 a_32668_n16916 0.285629f
C8737 a_44340_n3140 a_44452_n4328 0.026657f
C8738 a_23564_n17700 a_28076_n17349 0.028933f
C8739 a_37732_n20008 VDD 0.213126f
C8740 a_27572_860 a_28132_376 0.302602f
C8741 a_22444_n5156 a_23324_n7420 0.010366f
C8742 a_27988_n20388 a_28212_n20388 0.145671f
C8743 a_44788_n18820 a_45236_n18820 0.013276f
C8744 a_26271_n1400 VDD 0.572345f
C8745 a_43868_n20485 a_43780_n20388 0.285629f
C8746 a_45572_n9032 a_45660_n9076 0.285629f
C8747 a_46916_n9032 a_47364_n9032 0.013276f
C8748 a_28435_n10599 a_31961_n11340 0.013209f
C8749 a_44452_n10600 a_44092_n10644 0.086635f
C8750 a_43885_n452 a_43556_n661 0.014057f
C8751 a_21604_n8548 VDD 1.87917f
C8752 a_38268_n12212 a_38716_n12212 0.012882f
C8753 a_27281_n16854 a_27404_n14990 0.057877f
C8754 a_42660_n12168 a_42748_n12212 0.285629f
C8755 a_42100_n10980 VDD 0.205948f
C8756 a_32020_n2276 a_32432_n2689 0.536965f
C8757 a_38180_n15304 a_38628_n15304 0.013276f
C8758 a_40652_n1572 a_45572_n1192 0.049391f
C8759 a_43644_n705 a_43556_n661 0.49451f
C8760 a_34708_n17252 VDD 0.205948f
C8761 a_39972_n4328 a_40420_n4328 0.013276f
C8762 a_21792_n7464 a_21604_n5067 0.010233f
C8763 a_43644_n705 a_46243_769 0.037917f
C8764 a_40652_n1572 a_45212_332 0.029659f
C8765 a_44116_n5896 a_43756_n5940 0.086742f
C8766 a_33116_n18484 a_33564_n18484 0.012882f
C8767 a_42748_n7508 CLK 0.012909f
C8768 a_23844_n20008 a_23484_n20052 0.087066f
C8769 a_45212_n1669 VDD 0.316945f
C8770 a_40060_n9076 a_40172_n9509 0.026339f
C8771 a_44788_n4708 VDD 0.22479f
C8772 a_24965_n9860 a_23619_n12996 0.062527f
C8773 a_37732_n9032 VDD 0.213395f
C8774 a_47812_n12168 a_47452_n12212 0.086635f
C8775 a_40956_n13780 a_41404_n13780 0.012882f
C8776 a_31664_n13292 a_32413_n14564 0.063664f
C8777 a_21604_n708 a_22918_n2020 0.04208f
C8778 a_23912_n15216 VDD 0.3812f
C8779 a_41988_n2760 a_42436_n2760 0.013276f
C8780 a_22588_n18484 VDD 0.296789f
C8781 a_39056_820 a_38996_n408 0.032796f
C8782 a_23564_n17700 a_23844_n18440 0.038522f
C8783 a_42748_n16916 a_43196_n16916 0.012882f
C8784 a_34908_n16916 a_34796_n17349 0.026339f
C8785 a_39056_820 a_39544_420 0.08126f
C8786 a_47676_n20485 VDD 0.361497f
C8787 a_40420_n18440 a_40060_n18484 0.087066f
C8788 a_23887_n5156 a_24752_n8292 0.01296f
C8789 a_23479_n5156 a_26643_n8292 0.039375f
C8790 a_30340_n20008 a_30788_n20008 0.013276f
C8791 a_40532_n5896 VDD 0.207033f
C8792 a_25724_n14564 a_25132_n16432 0.117874f
C8793 a_30604_n11029 a_30296_n10980 0.934191f
C8794 a_47900_n9076 VDD 0.335152f
C8795 a_43644_n12212 a_43532_n12645 0.026339f
C8796 a_42300_n12212 VDD 0.315469f
C8797 a_37372_n13780 a_37484_n14213 0.026339f
C8798 a_29444_n708 a_29519_n1976 0.030366f
C8799 a_23404_816 a_25627_n452 0.041731f
C8800 a_42212_n15304 VDD 0.206217f
C8801 a_22140_n15781 a_22588_n15781 0.012552f
C8802 a_40652_n1572 a_41204_n1572 0.031385f
C8803 a_37284_n18440 VDD 0.231657f
C8804 a_27988_n4328 a_27597_n8292 0.014515f
C8805 a_22544_n4690 a_23887_n5156 0.031509f
C8806 a_41852_n16916 a_41740_n17349 0.026339f
C8807 a_47197_908 a_47924_376 0.168987f
C8808 a_36252_n18484 a_36140_n18917 0.026339f
C8809 a_45572_n18440 a_45660_n18484 0.285629f
C8810 a_46916_n18440 a_47364_n18440 0.013276f
C8811 a_30320_n6636 a_30740_n7464 0.097906f
C8812 a_30215_n6265 a_30111_n6221 0.277491f
C8813 a_42636_n7941 a_42996_n7844 0.087066f
C8814 a_27597_n8292 a_27485_n8500 0.026175f
C8815 a_24573_n6724 VDD 0.828867f
C8816 a_42636_n11077 a_43084_n11077 0.012882f
C8817 a_37036_n9509 VDD 0.33541f
C8818 a_30428_n12645 VDD 0.336455f
C8819 a_21916_n1975 a_26271_n1400 0.021843f
C8820 a_33452_n14213 a_33900_n14213 0.012882f
C8821 a_46556_n13780 a_46668_n14213 0.026339f
C8822 a_22948_n15684 VDD 0.207647f
C8823 a_27988_n4328 a_24492_n5156 0.074089f
C8824 a_26383_n2968 a_27337_n3140 0.020392f
C8825 a_25759_n3544 a_25600_n5895 0.019196f
C8826 a_23004_n2332 a_22820_n2804 0.075869f
C8827 a_21692_2431 a_28836_376 0.484278f
C8828 a_47900_n18484 VDD 0.335152f
C8829 a_29868_n17349 a_29780_n17252 0.285629f
C8830 a_40172_n17349 a_40620_n17349 0.012001f
C8831 a_46108_n4372 a_46220_n4805 0.026339f
C8832 a_47564_n6373 a_48012_n6373 0.012882f
C8833 a_43196_n18484 a_43084_n18917 0.026339f
C8834 a_22220_n9860 a_22264_n8988 0.131972f
C8835 a_42636_n6373 a_42548_n6276 0.285629f
C8836 a_44004_n20008 a_44452_n20008 0.013276f
C8837 a_40420_n20008 a_40508_n20052 0.285629f
C8838 a_28583_n3140 VDD 0.969759f
C8839 a_47116_n9509 a_47028_n9412 0.285629f
C8840 a_39188_n9412 a_39636_n9412 0.013276f
C8841 a_41204_n6276 VDD 0.227793f
C8842 a_45772_n11077 a_45684_n10980 0.285629f
C8843 a_37859_377 OUT[3] 0.139636f
C8844 a_43444_n9412 VDD 0.208665f
C8845 a_39500_n12645 a_39860_n12548 0.086742f
C8846 a_25132_n16432 a_25237_n13735 0.085656f
C8847 a_34932_n12548 VDD 0.209521f
C8848 a_35692_n14213 a_36052_n14116 0.087066f
C8849 a_35156_n15684 VDD 0.205948f
C8850 a_39724_n15781 a_39636_n15684 0.285629f
C8851 a_43084_n18917 VDD 0.313885f
C8852 a_40620_n17349 a_41204_n17252 0.016748f
C8853 a_23479_n5156 a_22264_n5852 0.250124f
C8854 a_41740_n4805 a_42188_n4805 0.012882f
C8855 a_46132_n4 a_46580_n4 0.013276f
C8856 a_23887_n5156 a_22016_n5825 0.04034f
C8857 a_25612_n18917 a_25972_n18820 0.087066f
C8858 a_38828_n18917 a_39276_n18917 0.012882f
C8859 a_46020_n20008 a_45660_n20052 0.086905f
C8860 a_39860_n7844 a_39972_n9032 0.026657f
C8861 XRST VSS 1.78628f
C8862 CLK VSS 9.525361f
C8863 EOC VSS 2.585921f
C8864 OUT[3] VSS 2.873034f
C8865 OUT[5] VSS 2.966969f
C8866 OUT[4] VSS 3.021139f
C8867 OUT[2] VSS 3.533625f
C8868 OUT[1] VSS 3.204847f
C8869 OUT[0] VSS 3.00522f
C8870 VIN VSS 1.35571f
C8871 VDD VSS 2.178174p
C8872 m3_n14480_n19265 VSS 4.74218f $ **FLOATING
C8873 m3_n14480_n16270 VSS 4.76818f $ **FLOATING
C8874 m3_n14480_n7750 VSS 4.704491f $ **FLOATING
C8875 m3_n14480_n4280 VSS 4.83805f $ **FLOATING
C8876 m3_n14480_n1270 VSS 4.73156f $ **FLOATING
C8877 a_47588_n20388 VSS 0.490237f
C8878 a_47140_n20388 VSS 0.478695f
C8879 a_46692_n20388 VSS 0.476546f
C8880 a_46244_n20388 VSS 0.475131f
C8881 a_45796_n20388 VSS 0.475131f
C8882 a_45348_n20388 VSS 0.475131f
C8883 a_44900_n20388 VSS 0.475131f
C8884 a_44452_n20388 VSS 0.487185f
C8885 a_43780_n20388 VSS 0.47896f
C8886 a_43332_n20388 VSS 0.476841f
C8887 a_42884_n20388 VSS 0.478828f
C8888 a_42436_n20388 VSS 0.479282f
C8889 a_41988_n20388 VSS 0.483976f
C8890 a_41540_n20388 VSS 0.510394f
C8891 a_41092_n20388 VSS 0.48209f
C8892 a_40644_n20388 VSS 0.491952f
C8893 a_39972_n20388 VSS 0.481297f
C8894 a_39524_n20388 VSS 0.475131f
C8895 a_39076_n20388 VSS 0.475131f
C8896 a_38628_n20388 VSS 0.475131f
C8897 a_38180_n20388 VSS 0.475131f
C8898 a_37732_n20388 VSS 0.475131f
C8899 a_37284_n20388 VSS 0.475131f
C8900 a_36836_n20388 VSS 0.487185f
C8901 a_36164_n20388 VSS 0.482371f
C8902 a_35716_n20388 VSS 0.480387f
C8903 a_35268_n20388 VSS 0.483211f
C8904 a_34820_n20388 VSS 0.518264f
C8905 a_34372_n20388 VSS 0.482683f
C8906 a_33924_n20388 VSS 0.480282f
C8907 a_33476_n20388 VSS 0.478512f
C8908 a_33028_n20388 VSS 0.488137f
C8909 a_32356_n20388 VSS 0.47896f
C8910 a_31908_n20388 VSS 0.475131f
C8911 a_31460_n20388 VSS 0.475131f
C8912 a_31012_n20388 VSS 0.475131f
C8913 a_30564_n20388 VSS 0.475131f
C8914 a_30116_n20388 VSS 0.475131f
C8915 a_29668_n20388 VSS 0.477348f
C8916 a_29220_n20388 VSS 0.496784f
C8917 a_28212_n20388 VSS 0.520474f
C8918 a_26756_n20388 VSS 0.488033f
C8919 a_26308_n20388 VSS 0.482148f
C8920 a_25860_n20388 VSS 0.480486f
C8921 a_25412_n20388 VSS 0.496661f
C8922 a_24516_n20388 VSS 0.495492f
C8923 a_47676_n20485 VSS 0.316718f
C8924 a_47228_n20485 VSS 0.29049f
C8925 a_46780_n20485 VSS 0.288809f
C8926 a_46332_n20485 VSS 0.2861f
C8927 a_45884_n20485 VSS 0.2861f
C8928 a_45436_n20485 VSS 0.2861f
C8929 a_44988_n20485 VSS 0.286193f
C8930 a_44540_n20485 VSS 0.284916f
C8931 a_43868_n20485 VSS 0.291256f
C8932 a_43420_n20485 VSS 0.287144f
C8933 a_42972_n20485 VSS 0.289911f
C8934 a_42524_n20485 VSS 0.291802f
C8935 a_42076_n20485 VSS 0.294175f
C8936 a_41628_n20485 VSS 0.333737f
C8937 a_41180_n20485 VSS 0.295027f
C8938 a_40732_n20485 VSS 0.295661f
C8939 a_40060_n20485 VSS 0.289403f
C8940 a_39612_n20485 VSS 0.281201f
C8941 a_39164_n20485 VSS 0.281201f
C8942 a_38716_n20485 VSS 0.281201f
C8943 a_38268_n20485 VSS 0.281201f
C8944 a_37820_n20485 VSS 0.281201f
C8945 a_37372_n20485 VSS 0.281201f
C8946 a_36924_n20485 VSS 0.289828f
C8947 a_36252_n20485 VSS 0.289734f
C8948 a_35804_n20485 VSS 0.286416f
C8949 a_35356_n20485 VSS 0.288686f
C8950 a_34908_n20485 VSS 0.314287f
C8951 a_34460_n20485 VSS 0.291084f
C8952 a_34012_n20485 VSS 0.2875f
C8953 a_33564_n20485 VSS 0.285361f
C8954 a_33116_n20485 VSS 0.286963f
C8955 a_32444_n20485 VSS 0.291173f
C8956 a_31996_n20485 VSS 0.286096f
C8957 a_31548_n20485 VSS 0.286096f
C8958 a_31100_n20485 VSS 0.286096f
C8959 a_30652_n20485 VSS 0.286096f
C8960 a_30204_n20485 VSS 0.286096f
C8961 a_29756_n20485 VSS 0.28766f
C8962 a_29308_n20485 VSS 0.294389f
C8963 a_28300_n20485 VSS 0.278985f
C8964 a_27540_n20747 VSS 0.434732f
C8965 a_26844_n20485 VSS 0.255089f
C8966 a_26396_n20485 VSS 0.29205f
C8967 a_25948_n20485 VSS 0.289078f
C8968 a_25500_n20485 VSS 0.292669f
C8969 a_24604_n20485 VSS 0.274557f
C8970 a_47900_n20052 VSS 0.305877f
C8971 a_47452_n20052 VSS 0.298988f
C8972 a_47004_n20052 VSS 0.296253f
C8973 a_46556_n20052 VSS 0.292631f
C8974 a_46108_n20052 VSS 0.290961f
C8975 a_45660_n20052 VSS 0.290961f
C8976 a_45212_n20052 VSS 0.29414f
C8977 a_47812_n20008 VSS 0.483823f
C8978 a_47364_n20008 VSS 0.46949f
C8979 a_46916_n20008 VSS 0.46798f
C8980 a_46468_n20008 VSS 0.461248f
C8981 a_46020_n20008 VSS 0.461248f
C8982 a_45572_n20008 VSS 0.461248f
C8983 a_45124_n20008 VSS 0.473068f
C8984 a_44540_n20052 VSS 0.287724f
C8985 a_44092_n20052 VSS 0.292638f
C8986 a_43644_n20052 VSS 0.289222f
C8987 a_43196_n20052 VSS 0.292271f
C8988 a_42748_n20052 VSS 0.29381f
C8989 a_42300_n20052 VSS 0.294653f
C8990 a_41852_n20052 VSS 0.305778f
C8991 a_41404_n20052 VSS 0.313702f
C8992 a_40956_n20052 VSS 0.296362f
C8993 a_40508_n20052 VSS 0.294065f
C8994 a_40060_n20052 VSS 0.285485f
C8995 a_39612_n20052 VSS 0.28236f
C8996 a_39164_n20052 VSS 0.28236f
C8997 a_38716_n20052 VSS 0.28236f
C8998 a_38268_n20052 VSS 0.28236f
C8999 a_37820_n20052 VSS 0.28236f
C9000 a_37372_n20052 VSS 0.285861f
C9001 a_44452_n20008 VSS 0.470565f
C9002 a_44004_n20008 VSS 0.45666f
C9003 a_43556_n20008 VSS 0.45666f
C9004 a_43108_n20008 VSS 0.459647f
C9005 a_42660_n20008 VSS 0.461258f
C9006 a_42212_n20008 VSS 0.462696f
C9007 a_41764_n20008 VSS 0.485271f
C9008 a_41316_n20008 VSS 0.465969f
C9009 a_40868_n20008 VSS 0.477382f
C9010 a_40420_n20008 VSS 0.461802f
C9011 a_39972_n20008 VSS 0.460237f
C9012 a_39524_n20008 VSS 0.4579f
C9013 a_39076_n20008 VSS 0.4579f
C9014 a_38628_n20008 VSS 0.4579f
C9015 a_38180_n20008 VSS 0.4579f
C9016 a_37732_n20008 VSS 0.4579f
C9017 a_37284_n20008 VSS 0.46986f
C9018 a_36700_n20052 VSS 0.294796f
C9019 a_36252_n20052 VSS 0.289297f
C9020 a_35804_n20052 VSS 0.287575f
C9021 a_35356_n20052 VSS 0.289845f
C9022 a_34908_n20052 VSS 0.315438f
C9023 a_34460_n20052 VSS 0.292218f
C9024 a_34012_n20052 VSS 0.288659f
C9025 a_33564_n20052 VSS 0.28652f
C9026 a_33116_n20052 VSS 0.284407f
C9027 a_32668_n20052 VSS 0.289158f
C9028 a_32220_n20052 VSS 0.289222f
C9029 a_31772_n20052 VSS 0.289222f
C9030 a_31324_n20052 VSS 0.289222f
C9031 a_30876_n20052 VSS 0.289222f
C9032 a_30428_n20052 VSS 0.289222f
C9033 a_29980_n20052 VSS 0.289222f
C9034 a_29532_n20052 VSS 0.295928f
C9035 a_36612_n20008 VSS 0.471561f
C9036 a_36164_n20008 VSS 0.460071f
C9037 a_35716_n20008 VSS 0.461917f
C9038 a_35268_n20008 VSS 0.464741f
C9039 a_34820_n20008 VSS 0.50076f
C9040 a_34372_n20008 VSS 0.464212f
C9041 a_33924_n20008 VSS 0.461811f
C9042 a_33476_n20008 VSS 0.460042f
C9043 a_33028_n20008 VSS 0.472504f
C9044 a_32580_n20008 VSS 0.457943f
C9045 a_32132_n20008 VSS 0.4579f
C9046 a_31684_n20008 VSS 0.4579f
C9047 a_31236_n20008 VSS 0.4579f
C9048 a_30788_n20008 VSS 0.4579f
C9049 a_30340_n20008 VSS 0.4579f
C9050 a_29892_n20008 VSS 0.458024f
C9051 a_29444_n20008 VSS 0.473009f
C9052 a_28860_n20052 VSS 0.300426f
C9053 a_28412_n20052 VSS 0.298078f
C9054 a_27964_n20052 VSS 0.326219f
C9055 a_27516_n20052 VSS 0.293915f
C9056 a_27068_n20052 VSS 0.294625f
C9057 a_26620_n20052 VSS 0.292876f
C9058 a_26172_n20052 VSS 0.289827f
C9059 a_25724_n20052 VSS 0.289229f
C9060 a_25276_n20052 VSS 0.289321f
C9061 a_24828_n20052 VSS 0.289066f
C9062 a_24380_n20052 VSS 0.289356f
C9063 a_23932_n20052 VSS 0.28236f
C9064 a_23484_n20052 VSS 0.285163f
C9065 a_23036_n20052 VSS 0.28236f
C9066 a_22588_n20052 VSS 0.28236f
C9067 a_22140_n20052 VSS 0.28236f
C9068 a_21692_n20052 VSS 0.295089f
C9069 a_28772_n20008 VSS 0.477882f
C9070 a_28324_n20008 VSS 0.466575f
C9071 a_27876_n20008 VSS 0.481423f
C9072 a_27428_n20008 VSS 0.463608f
C9073 a_26980_n20008 VSS 0.461473f
C9074 a_26532_n20008 VSS 0.46098f
C9075 a_26084_n20008 VSS 0.45666f
C9076 a_25636_n20008 VSS 0.45666f
C9077 a_25188_n20008 VSS 0.471552f
C9078 a_24740_n20008 VSS 0.440291f
C9079 a_24292_n20008 VSS 0.440291f
C9080 a_23844_n20008 VSS 0.440291f
C9081 a_23396_n20008 VSS 0.440291f
C9082 a_22948_n20008 VSS 0.440291f
C9083 a_22500_n20008 VSS 0.440291f
C9084 a_22052_n20008 VSS 0.440291f
C9085 a_21604_n20008 VSS 0.468317f
C9086 a_47924_n18820 VSS 0.475688f
C9087 a_47476_n18820 VSS 0.461842f
C9088 a_47028_n18820 VSS 0.460159f
C9089 a_46580_n18820 VSS 0.45746f
C9090 a_46132_n18820 VSS 0.45695f
C9091 a_45684_n18820 VSS 0.45695f
C9092 a_45236_n18820 VSS 0.45695f
C9093 a_44788_n18820 VSS 0.472938f
C9094 a_44340_n18820 VSS 0.459328f
C9095 a_43892_n18820 VSS 0.458189f
C9096 a_43444_n18820 VSS 0.458947f
C9097 a_42996_n18820 VSS 0.461509f
C9098 a_42548_n18820 VSS 0.463309f
C9099 a_42100_n18820 VSS 0.466069f
C9100 a_41652_n18820 VSS 0.499854f
C9101 a_41204_n18820 VSS 0.477949f
C9102 a_40532_n18820 VSS 0.475145f
C9103 a_40084_n18820 VSS 0.460833f
C9104 a_39636_n18820 VSS 0.45801f
C9105 a_39188_n18820 VSS 0.45801f
C9106 a_38740_n18820 VSS 0.45801f
C9107 a_38292_n18820 VSS 0.45801f
C9108 a_37844_n18820 VSS 0.45801f
C9109 a_37396_n18820 VSS 0.45801f
C9110 a_36948_n18820 VSS 0.472902f
C9111 a_36500_n18820 VSS 0.461296f
C9112 a_36052_n18820 VSS 0.463085f
C9113 a_35604_n18820 VSS 0.465108f
C9114 a_35156_n18820 VSS 0.468594f
C9115 a_34708_n18820 VSS 0.492113f
C9116 a_34260_n18820 VSS 0.466082f
C9117 a_33812_n18820 VSS 0.463929f
C9118 a_33364_n18820 VSS 0.474293f
C9119 a_32692_n18820 VSS 0.471958f
C9120 a_32244_n18820 VSS 0.45695f
C9121 a_31796_n18820 VSS 0.45695f
C9122 a_31348_n18820 VSS 0.45695f
C9123 a_30900_n18820 VSS 0.45695f
C9124 a_30452_n18820 VSS 0.45695f
C9125 a_30004_n18820 VSS 0.45695f
C9126 a_29556_n18820 VSS 0.459785f
C9127 a_29108_n18820 VSS 0.477292f
C9128 a_28660_n18820 VSS 0.46593f
C9129 a_28212_n18820 VSS 0.480167f
C9130 a_27764_n18820 VSS 0.47113f
C9131 a_27316_n18820 VSS 0.465358f
C9132 a_26868_n18820 VSS 0.462258f
C9133 a_26420_n18820 VSS 0.460873f
C9134 a_25972_n18820 VSS 0.458189f
C9135 a_25524_n18820 VSS 0.472692f
C9136 a_24740_n18820 VSS 0.442147f
C9137 a_24292_n18820 VSS 0.438283f
C9138 a_23844_n18820 VSS 0.438283f
C9139 a_23396_n18820 VSS 0.438283f
C9140 a_22948_n18820 VSS 0.438283f
C9141 a_22500_n18820 VSS 0.438283f
C9142 a_22052_n18820 VSS 0.438283f
C9143 a_21604_n18820 VSS 0.466401f
C9144 a_48012_n18917 VSS 0.321039f
C9145 a_47564_n18917 VSS 0.290098f
C9146 a_47116_n18917 VSS 0.288045f
C9147 a_46668_n18917 VSS 0.28552f
C9148 a_46220_n18917 VSS 0.284099f
C9149 a_45772_n18917 VSS 0.284099f
C9150 a_45324_n18917 VSS 0.284099f
C9151 a_44876_n18917 VSS 0.285753f
C9152 a_44428_n18917 VSS 0.284269f
C9153 a_43980_n18917 VSS 0.284258f
C9154 a_43532_n18917 VSS 0.284258f
C9155 a_43084_n18917 VSS 0.287629f
C9156 a_42636_n18917 VSS 0.289343f
C9157 a_42188_n18917 VSS 0.290362f
C9158 a_41740_n18917 VSS 0.314383f
C9159 a_41292_n18917 VSS 0.298098f
C9160 a_40620_n18917 VSS 0.294742f
C9161 a_40172_n18917 VSS 0.291042f
C9162 a_39724_n18917 VSS 0.284188f
C9163 a_39276_n18917 VSS 0.284099f
C9164 a_38828_n18917 VSS 0.284099f
C9165 a_38380_n18917 VSS 0.284099f
C9166 a_37932_n18917 VSS 0.284099f
C9167 a_37484_n18917 VSS 0.284099f
C9168 a_37036_n18917 VSS 0.285753f
C9169 a_36588_n18917 VSS 0.28553f
C9170 a_36140_n18917 VSS 0.288087f
C9171 a_35692_n18917 VSS 0.29002f
C9172 a_35244_n18917 VSS 0.292499f
C9173 a_34796_n18917 VSS 0.331502f
C9174 a_34348_n18917 VSS 0.292838f
C9175 a_33900_n18917 VSS 0.289962f
C9176 a_33452_n18917 VSS 0.291503f
C9177 a_32780_n18917 VSS 0.291094f
C9178 a_32332_n18917 VSS 0.289297f
C9179 a_31884_n18917 VSS 0.285816f
C9180 a_31436_n18917 VSS 0.285816f
C9181 a_30988_n18917 VSS 0.285812f
C9182 a_30540_n18917 VSS 0.285812f
C9183 a_30092_n18917 VSS 0.285812f
C9184 a_29644_n18917 VSS 0.28855f
C9185 a_29196_n18917 VSS 0.293103f
C9186 a_28748_n18917 VSS 0.294943f
C9187 a_28300_n18917 VSS 0.2987f
C9188 a_27852_n18917 VSS 0.320332f
C9189 a_27404_n18917 VSS 0.296104f
C9190 a_26956_n18917 VSS 0.293549f
C9191 a_26508_n18917 VSS 0.291666f
C9192 a_26060_n18917 VSS 0.285899f
C9193 a_25612_n18917 VSS 0.289629f
C9194 a_24828_n18917 VSS 0.269581f
C9195 a_24380_n18917 VSS 0.281201f
C9196 a_23932_n18917 VSS 0.281201f
C9197 a_23484_n18917 VSS 0.281201f
C9198 a_23036_n18917 VSS 0.281201f
C9199 a_22588_n18917 VSS 0.281201f
C9200 a_22140_n18917 VSS 0.281201f
C9201 a_21692_n18917 VSS 0.291339f
C9202 a_47900_n18484 VSS 0.300977f
C9203 a_47452_n18484 VSS 0.294024f
C9204 a_47004_n18484 VSS 0.29129f
C9205 a_46556_n18484 VSS 0.287668f
C9206 a_46108_n18484 VSS 0.285997f
C9207 a_45660_n18484 VSS 0.285997f
C9208 a_45212_n18484 VSS 0.289177f
C9209 a_47812_n18440 VSS 0.483823f
C9210 a_47364_n18440 VSS 0.46949f
C9211 a_46916_n18440 VSS 0.46798f
C9212 a_46468_n18440 VSS 0.461248f
C9213 a_46020_n18440 VSS 0.461248f
C9214 a_45572_n18440 VSS 0.461248f
C9215 a_45124_n18440 VSS 0.473068f
C9216 a_44540_n18484 VSS 0.289463f
C9217 a_44092_n18484 VSS 0.287579f
C9218 a_43644_n18484 VSS 0.284099f
C9219 a_43196_n18484 VSS 0.287148f
C9220 a_42748_n18484 VSS 0.288687f
C9221 a_42300_n18484 VSS 0.28953f
C9222 a_41852_n18484 VSS 0.300321f
C9223 a_41404_n18484 VSS 0.308618f
C9224 a_40956_n18484 VSS 0.292892f
C9225 a_40508_n18484 VSS 0.289019f
C9226 a_40060_n18484 VSS 0.287384f
C9227 a_39612_n18484 VSS 0.284258f
C9228 a_39164_n18484 VSS 0.284258f
C9229 a_38716_n18484 VSS 0.284258f
C9230 a_38268_n18484 VSS 0.284258f
C9231 a_37820_n18484 VSS 0.284258f
C9232 a_37372_n18484 VSS 0.287759f
C9233 a_44452_n18440 VSS 0.470565f
C9234 a_44004_n18440 VSS 0.45666f
C9235 a_43556_n18440 VSS 0.45666f
C9236 a_43108_n18440 VSS 0.459647f
C9237 a_42660_n18440 VSS 0.461258f
C9238 a_42212_n18440 VSS 0.462696f
C9239 a_41764_n18440 VSS 0.485271f
C9240 a_41316_n18440 VSS 0.465969f
C9241 a_40868_n18440 VSS 0.477382f
C9242 a_40420_n18440 VSS 0.461802f
C9243 a_39972_n18440 VSS 0.460237f
C9244 a_39524_n18440 VSS 0.4579f
C9245 a_39076_n18440 VSS 0.4579f
C9246 a_38628_n18440 VSS 0.4579f
C9247 a_38180_n18440 VSS 0.4579f
C9248 a_37732_n18440 VSS 0.4579f
C9249 a_37284_n18440 VSS 0.46986f
C9250 a_36700_n18484 VSS 0.289581f
C9251 a_36252_n18484 VSS 0.291036f
C9252 a_35804_n18484 VSS 0.289314f
C9253 a_35356_n18484 VSS 0.291585f
C9254 a_34908_n18484 VSS 0.318139f
C9255 a_34460_n18484 VSS 0.293957f
C9256 a_34012_n18484 VSS 0.290398f
C9257 a_33564_n18484 VSS 0.288259f
C9258 a_33116_n18484 VSS 0.2878f
C9259 a_32668_n18484 VSS 0.284269f
C9260 a_32220_n18484 VSS 0.284258f
C9261 a_31772_n18484 VSS 0.284258f
C9262 a_31324_n18484 VSS 0.284258f
C9263 a_30876_n18484 VSS 0.284258f
C9264 a_30428_n18484 VSS 0.284258f
C9265 a_29980_n18484 VSS 0.284258f
C9266 a_29532_n18484 VSS 0.29152f
C9267 a_36612_n18440 VSS 0.471561f
C9268 a_36164_n18440 VSS 0.460071f
C9269 a_35716_n18440 VSS 0.461917f
C9270 a_35268_n18440 VSS 0.464741f
C9271 a_34820_n18440 VSS 0.50076f
C9272 a_34372_n18440 VSS 0.464212f
C9273 a_33924_n18440 VSS 0.461811f
C9274 a_33476_n18440 VSS 0.460042f
C9275 a_33028_n18440 VSS 0.472504f
C9276 a_32580_n18440 VSS 0.45666f
C9277 a_32132_n18440 VSS 0.45666f
C9278 a_31684_n18440 VSS 0.45666f
C9279 a_31236_n18440 VSS 0.45666f
C9280 a_30788_n18440 VSS 0.45666f
C9281 a_30340_n18440 VSS 0.45666f
C9282 a_29892_n18440 VSS 0.458135f
C9283 a_29444_n18440 VSS 0.478813f
C9284 a_28524_n18484 VSS 0.278515f
C9285 a_28076_n18484 VSS 0.327517f
C9286 a_27628_n18484 VSS 0.29669f
C9287 a_27180_n18484 VSS 0.295009f
C9288 a_26172_n18484 VSS 0.25765f
C9289 a_25724_n18484 VSS 0.288447f
C9290 a_25276_n18484 VSS 0.289231f
C9291 a_24828_n18484 VSS 0.284681f
C9292 a_24380_n18484 VSS 0.281201f
C9293 a_23932_n18484 VSS 0.281201f
C9294 a_23484_n18484 VSS 0.281201f
C9295 a_23036_n18484 VSS 0.281201f
C9296 a_22588_n18484 VSS 0.281201f
C9297 a_22140_n18484 VSS 0.281201f
C9298 a_21692_n18484 VSS 0.291339f
C9299 a_28436_n18440 VSS 0.456176f
C9300 a_27988_n18440 VSS 0.486902f
C9301 a_27540_n18440 VSS 0.481247f
C9302 a_27092_n18440 VSS 0.495721f
C9303 a_26084_n18440 VSS 0.484415f
C9304 a_25636_n18440 VSS 0.477732f
C9305 a_25188_n18440 VSS 0.481183f
C9306 a_24740_n18440 VSS 0.46996f
C9307 a_24292_n18440 VSS 0.472379f
C9308 a_23844_n18440 VSS 0.450965f
C9309 a_23396_n18440 VSS 0.451147f
C9310 a_22948_n18440 VSS 0.451008f
C9311 a_22500_n18440 VSS 0.451008f
C9312 a_22052_n18440 VSS 0.451008f
C9313 a_21604_n18440 VSS 0.479265f
C9314 a_47924_n17252 VSS 0.474295f
C9315 a_47476_n17252 VSS 0.461553f
C9316 a_47028_n17252 VSS 0.45987f
C9317 a_46580_n17252 VSS 0.457171f
C9318 a_46132_n17252 VSS 0.45666f
C9319 a_45684_n17252 VSS 0.45666f
C9320 a_45236_n17252 VSS 0.45666f
C9321 a_44788_n17252 VSS 0.471552f
C9322 a_44340_n17252 VSS 0.457943f
C9323 a_43892_n17252 VSS 0.4579f
C9324 a_43444_n17252 VSS 0.458658f
C9325 a_42996_n17252 VSS 0.46122f
C9326 a_42548_n17252 VSS 0.463019f
C9327 a_42100_n17252 VSS 0.46578f
C9328 a_41652_n17252 VSS 0.499395f
C9329 a_41204_n17252 VSS 0.47766f
C9330 a_40532_n17252 VSS 0.474856f
C9331 a_40084_n17252 VSS 0.459483f
C9332 a_39636_n17252 VSS 0.45666f
C9333 a_39188_n17252 VSS 0.45666f
C9334 a_38740_n17252 VSS 0.45666f
C9335 a_38292_n17252 VSS 0.45666f
C9336 a_37844_n17252 VSS 0.45666f
C9337 a_37396_n17252 VSS 0.45666f
C9338 a_36948_n17252 VSS 0.471552f
C9339 a_36500_n17252 VSS 0.459903f
C9340 a_36052_n17252 VSS 0.461699f
C9341 a_35604_n17252 VSS 0.463723f
C9342 a_35156_n17252 VSS 0.467208f
C9343 a_34708_n17252 VSS 0.490181f
C9344 a_34260_n17252 VSS 0.464697f
C9345 a_33812_n17252 VSS 0.462544f
C9346 a_33364_n17252 VSS 0.477263f
C9347 a_32468_n17252 VSS 0.47335f
C9348 a_32020_n17252 VSS 0.466435f
C9349 a_31572_n17252 VSS 0.466435f
C9350 a_31124_n17252 VSS 0.457242f
C9351 a_30676_n17252 VSS 0.457242f
C9352 a_30228_n17252 VSS 0.457242f
C9353 a_29780_n17252 VSS 0.458471f
C9354 a_29332_n17252 VSS 0.460746f
C9355 a_28884_n17252 VSS 0.475356f
C9356 a_28436_n17252 VSS 0.446297f
C9357 a_27988_n17252 VSS 0.506649f
C9358 a_24516_n17252 VSS 0.494417f
C9359 a_48012_n17349 VSS 0.321039f
C9360 a_47564_n17349 VSS 0.290098f
C9361 a_47116_n17349 VSS 0.288045f
C9362 a_46668_n17349 VSS 0.28552f
C9363 a_46220_n17349 VSS 0.284099f
C9364 a_45772_n17349 VSS 0.284099f
C9365 a_45324_n17349 VSS 0.284099f
C9366 a_44876_n17349 VSS 0.285753f
C9367 a_44428_n17349 VSS 0.284269f
C9368 a_43980_n17349 VSS 0.284258f
C9369 a_43532_n17349 VSS 0.284258f
C9370 a_43084_n17349 VSS 0.287629f
C9371 a_42636_n17349 VSS 0.289343f
C9372 a_42188_n17349 VSS 0.290362f
C9373 a_41740_n17349 VSS 0.314383f
C9374 a_41292_n17349 VSS 0.298098f
C9375 a_40620_n17349 VSS 0.294742f
C9376 a_40172_n17349 VSS 0.291042f
C9377 a_39724_n17349 VSS 0.284188f
C9378 a_39276_n17349 VSS 0.284099f
C9379 a_38828_n17349 VSS 0.284099f
C9380 a_38380_n17349 VSS 0.284099f
C9381 a_37932_n17349 VSS 0.284099f
C9382 a_37484_n17349 VSS 0.284099f
C9383 a_37036_n17349 VSS 0.285753f
C9384 a_36588_n17349 VSS 0.28553f
C9385 a_36140_n17349 VSS 0.288095f
C9386 a_35692_n17349 VSS 0.290028f
C9387 a_35244_n17349 VSS 0.292503f
C9388 a_34796_n17349 VSS 0.331503f
C9389 a_34348_n17349 VSS 0.292842f
C9390 a_33900_n17349 VSS 0.289966f
C9391 a_33452_n17349 VSS 0.291912f
C9392 a_32556_n17349 VSS 0.271024f
C9393 a_32108_n17349 VSS 0.288936f
C9394 a_31660_n17349 VSS 0.288066f
C9395 a_31212_n17349 VSS 0.286908f
C9396 a_30764_n17349 VSS 0.283428f
C9397 a_30316_n17349 VSS 0.283686f
C9398 a_29868_n17349 VSS 0.285457f
C9399 a_29420_n17349 VSS 0.290874f
C9400 a_28972_n17349 VSS 0.291093f
C9401 a_28524_n17349 VSS 0.289885f
C9402 a_28076_n17349 VSS 0.321564f
C9403 a_24604_n17349 VSS 0.273552f
C9404 a_47900_n16916 VSS 0.300977f
C9405 a_47452_n16916 VSS 0.294024f
C9406 a_47004_n16916 VSS 0.29129f
C9407 a_46556_n16916 VSS 0.287668f
C9408 a_46108_n16916 VSS 0.285997f
C9409 a_45660_n16916 VSS 0.285997f
C9410 a_45212_n16916 VSS 0.289177f
C9411 a_47812_n16872 VSS 0.483823f
C9412 a_47364_n16872 VSS 0.46949f
C9413 a_46916_n16872 VSS 0.46798f
C9414 a_46468_n16872 VSS 0.461248f
C9415 a_46020_n16872 VSS 0.461248f
C9416 a_45572_n16872 VSS 0.461248f
C9417 a_45124_n16872 VSS 0.473068f
C9418 a_44540_n16916 VSS 0.289463f
C9419 a_44092_n16916 VSS 0.287579f
C9420 a_43644_n16916 VSS 0.284099f
C9421 a_43196_n16916 VSS 0.287148f
C9422 a_42748_n16916 VSS 0.288687f
C9423 a_42300_n16916 VSS 0.28953f
C9424 a_41852_n16916 VSS 0.300321f
C9425 a_41404_n16916 VSS 0.308618f
C9426 a_40956_n16916 VSS 0.292892f
C9427 a_40508_n16916 VSS 0.289019f
C9428 a_40060_n16916 VSS 0.287384f
C9429 a_39612_n16916 VSS 0.284258f
C9430 a_39164_n16916 VSS 0.284258f
C9431 a_38716_n16916 VSS 0.284258f
C9432 a_38268_n16916 VSS 0.284258f
C9433 a_37820_n16916 VSS 0.284258f
C9434 a_37372_n16916 VSS 0.287759f
C9435 a_44452_n16872 VSS 0.470565f
C9436 a_44004_n16872 VSS 0.45666f
C9437 a_43556_n16872 VSS 0.45666f
C9438 a_43108_n16872 VSS 0.459647f
C9439 a_42660_n16872 VSS 0.461258f
C9440 a_42212_n16872 VSS 0.462696f
C9441 a_41764_n16872 VSS 0.485271f
C9442 a_41316_n16872 VSS 0.465969f
C9443 a_40868_n16872 VSS 0.477382f
C9444 a_40420_n16872 VSS 0.461802f
C9445 a_39972_n16872 VSS 0.460237f
C9446 a_39524_n16872 VSS 0.4579f
C9447 a_39076_n16872 VSS 0.4579f
C9448 a_38628_n16872 VSS 0.4579f
C9449 a_38180_n16872 VSS 0.4579f
C9450 a_37732_n16872 VSS 0.4579f
C9451 a_37284_n16872 VSS 0.46986f
C9452 a_36700_n16916 VSS 0.289581f
C9453 a_36252_n16916 VSS 0.291904f
C9454 a_35804_n16916 VSS 0.292792f
C9455 a_35356_n16916 VSS 0.294629f
C9456 a_34908_n16916 VSS 0.319866f
C9457 a_34460_n16916 VSS 0.295657f
C9458 a_34012_n16916 VSS 0.292137f
C9459 a_33564_n16916 VSS 0.289275f
C9460 a_33116_n16916 VSS 0.286641f
C9461 a_32668_n16916 VSS 0.28294f
C9462 a_32220_n16916 VSS 0.28294f
C9463 a_31772_n16916 VSS 0.28294f
C9464 a_31324_n16916 VSS 0.28294f
C9465 a_30876_n16916 VSS 0.28294f
C9466 a_30428_n16916 VSS 0.2828f
C9467 a_36612_n16872 VSS 0.472912f
C9468 a_36164_n16872 VSS 0.468606f
C9469 a_35716_n16872 VSS 0.470452f
C9470 a_35268_n16872 VSS 0.469439f
C9471 a_34820_n16872 VSS 0.505933f
C9472 a_34372_n16872 VSS 0.468911f
C9473 a_33924_n16872 VSS 0.466509f
C9474 a_33476_n16872 VSS 0.459384f
C9475 a_33028_n16872 VSS 0.471846f
C9476 a_32580_n16872 VSS 0.469442f
C9477 a_32132_n16872 VSS 0.466262f
C9478 a_31684_n16872 VSS 0.462587f
C9479 a_31236_n16872 VSS 0.462587f
C9480 a_30788_n16872 VSS 0.462587f
C9481 a_30340_n16872 VSS 0.486556f
C9482 a_28636_n16916 VSS 0.248786f
C9483 a_25544_n16412 VSS 0.41419f
C9484 a_23932_n16916 VSS 0.239679f
C9485 a_23484_n16916 VSS 0.287202f
C9486 a_23036_n16916 VSS 0.285404f
C9487 a_22588_n16916 VSS 0.284099f
C9488 a_22140_n16916 VSS 0.284099f
C9489 a_21692_n16916 VSS 0.295068f
C9490 a_28548_n16872 VSS 0.501427f
C9491 a_23844_n16872 VSS 0.4772f
C9492 a_23396_n16872 VSS 0.476707f
C9493 a_22948_n16872 VSS 0.443639f
C9494 a_22500_n16872 VSS 0.443639f
C9495 a_22052_n16872 VSS 0.443639f
C9496 a_21604_n16872 VSS 0.471527f
C9497 a_47924_n15684 VSS 0.474295f
C9498 a_47476_n15684 VSS 0.461553f
C9499 a_47028_n15684 VSS 0.45987f
C9500 a_46580_n15684 VSS 0.457171f
C9501 a_46132_n15684 VSS 0.45666f
C9502 a_45684_n15684 VSS 0.45666f
C9503 a_45236_n15684 VSS 0.45666f
C9504 a_44788_n15684 VSS 0.471552f
C9505 a_44340_n15684 VSS 0.457943f
C9506 a_43892_n15684 VSS 0.4579f
C9507 a_43444_n15684 VSS 0.458658f
C9508 a_42996_n15684 VSS 0.46122f
C9509 a_42548_n15684 VSS 0.463019f
C9510 a_42100_n15684 VSS 0.46578f
C9511 a_41652_n15684 VSS 0.499395f
C9512 a_41204_n15684 VSS 0.47766f
C9513 a_40532_n15684 VSS 0.474856f
C9514 a_40084_n15684 VSS 0.459483f
C9515 a_39636_n15684 VSS 0.45666f
C9516 a_39188_n15684 VSS 0.45666f
C9517 a_38740_n15684 VSS 0.45666f
C9518 a_38292_n15684 VSS 0.45666f
C9519 a_37844_n15684 VSS 0.45666f
C9520 a_37396_n15684 VSS 0.45666f
C9521 a_36948_n15684 VSS 0.471552f
C9522 a_36500_n15684 VSS 0.459903f
C9523 a_36052_n15684 VSS 0.461732f
C9524 a_35604_n15684 VSS 0.463755f
C9525 a_35156_n15684 VSS 0.467225f
C9526 a_34708_n15684 VSS 0.490107f
C9527 a_34260_n15684 VSS 0.464713f
C9528 a_33812_n15684 VSS 0.46256f
C9529 a_33364_n15684 VSS 0.479083f
C9530 a_23564_n17700 VSS 2.06881f
C9531 a_48012_n15781 VSS 0.321039f
C9532 a_47564_n15781 VSS 0.290098f
C9533 a_47116_n15781 VSS 0.288045f
C9534 a_46668_n15781 VSS 0.28552f
C9535 a_46220_n15781 VSS 0.284099f
C9536 a_45772_n15781 VSS 0.284099f
C9537 a_45324_n15781 VSS 0.284099f
C9538 a_44876_n15781 VSS 0.285753f
C9539 a_44428_n15781 VSS 0.284269f
C9540 a_43980_n15781 VSS 0.284258f
C9541 a_43532_n15781 VSS 0.284258f
C9542 a_43084_n15781 VSS 0.287629f
C9543 a_42636_n15781 VSS 0.289343f
C9544 a_42188_n15781 VSS 0.290362f
C9545 a_41740_n15781 VSS 0.314383f
C9546 a_41292_n15781 VSS 0.298098f
C9547 a_40620_n15781 VSS 0.294742f
C9548 a_40172_n15781 VSS 0.291042f
C9549 a_39724_n15781 VSS 0.284188f
C9550 a_39276_n15781 VSS 0.284099f
C9551 a_38828_n15781 VSS 0.284099f
C9552 a_38380_n15781 VSS 0.284099f
C9553 a_37932_n15781 VSS 0.284099f
C9554 a_37484_n15781 VSS 0.284099f
C9555 a_37036_n15781 VSS 0.285753f
C9556 a_36588_n15781 VSS 0.283621f
C9557 a_36140_n15781 VSS 0.286189f
C9558 a_35692_n15781 VSS 0.288122f
C9559 a_35244_n15781 VSS 0.290601f
C9560 a_34796_n15781 VSS 0.328462f
C9561 a_34348_n15781 VSS 0.29094f
C9562 a_33900_n15781 VSS 0.288064f
C9563 a_33452_n15781 VSS 0.289986f
C9564 a_28568_n16066 VSS 0.715069f
C9565 a_27709_n16132 VSS 0.797929f
C9566 a_27085_n16132 VSS 0.771934f
C9567 a_23564_n20836 VSS 2.10484f
C9568 a_22948_n15684 VSS 0.448123f
C9569 a_22500_n15684 VSS 0.443639f
C9570 a_22052_n15684 VSS 0.443639f
C9571 a_21604_n15684 VSS 0.471527f
C9572 a_26755_n16132 VSS 0.636966f
C9573 a_24752_n16132 VSS 0.389616f
C9574 a_24088_n16087 VSS 0.414865f
C9575 a_23036_n15781 VSS 0.252822f
C9576 a_22588_n15781 VSS 0.285923f
C9577 a_22140_n15781 VSS 0.284099f
C9578 a_21692_n15781 VSS 0.293704f
C9579 a_47900_n15348 VSS 0.300977f
C9580 a_47452_n15348 VSS 0.294024f
C9581 a_47004_n15348 VSS 0.29129f
C9582 a_46556_n15348 VSS 0.287668f
C9583 a_46108_n15348 VSS 0.285997f
C9584 a_45660_n15348 VSS 0.285997f
C9585 a_45212_n15348 VSS 0.289177f
C9586 a_47812_n15304 VSS 0.483823f
C9587 a_47364_n15304 VSS 0.46949f
C9588 a_46916_n15304 VSS 0.46798f
C9589 a_46468_n15304 VSS 0.461248f
C9590 a_46020_n15304 VSS 0.461248f
C9591 a_45572_n15304 VSS 0.461248f
C9592 a_45124_n15304 VSS 0.473068f
C9593 a_44540_n15348 VSS 0.289463f
C9594 a_44092_n15348 VSS 0.287579f
C9595 a_43644_n15348 VSS 0.284099f
C9596 a_43196_n15348 VSS 0.287148f
C9597 a_42748_n15348 VSS 0.288687f
C9598 a_42300_n15348 VSS 0.28953f
C9599 a_41852_n15348 VSS 0.300321f
C9600 a_41404_n15348 VSS 0.308618f
C9601 a_40956_n15348 VSS 0.292892f
C9602 a_40508_n15348 VSS 0.289019f
C9603 a_40060_n15348 VSS 0.287384f
C9604 a_39612_n15348 VSS 0.284258f
C9605 a_39164_n15348 VSS 0.284258f
C9606 a_38716_n15348 VSS 0.284258f
C9607 a_38268_n15348 VSS 0.284258f
C9608 a_37820_n15348 VSS 0.284258f
C9609 a_37372_n15348 VSS 0.287991f
C9610 a_44452_n15304 VSS 0.470565f
C9611 a_44004_n15304 VSS 0.45666f
C9612 a_43556_n15304 VSS 0.45666f
C9613 a_43108_n15304 VSS 0.459647f
C9614 a_42660_n15304 VSS 0.461258f
C9615 a_42212_n15304 VSS 0.462696f
C9616 a_41764_n15304 VSS 0.485271f
C9617 a_41316_n15304 VSS 0.465969f
C9618 a_40868_n15304 VSS 0.477382f
C9619 a_40420_n15304 VSS 0.461802f
C9620 a_39972_n15304 VSS 0.460237f
C9621 a_39524_n15304 VSS 0.4579f
C9622 a_39076_n15304 VSS 0.4579f
C9623 a_38628_n15304 VSS 0.4579f
C9624 a_38180_n15304 VSS 0.4579f
C9625 a_37732_n15304 VSS 0.4579f
C9626 a_37284_n15304 VSS 0.472403f
C9627 a_36588_n15348 VSS 0.272289f
C9628 a_36140_n15348 VSS 0.28938f
C9629 a_35692_n15348 VSS 0.286963f
C9630 a_35244_n15348 VSS 0.289445f
C9631 a_34796_n15348 VSS 0.324566f
C9632 a_34348_n15348 VSS 0.288978f
C9633 a_33900_n15348 VSS 0.286289f
C9634 a_33452_n15348 VSS 0.284522f
C9635 a_33004_n15348 VSS 0.287924f
C9636 a_28212_n15303 VSS 0.011683f
C9637 a_27988_n20388 VSS 2.47608f
C9638 a_36500_n15304 VSS 0.45619f
C9639 a_36052_n15304 VSS 0.442083f
C9640 a_35604_n15304 VSS 0.444106f
C9641 a_35156_n15304 VSS 0.445882f
C9642 a_34708_n15304 VSS 0.468367f
C9643 a_34260_n15304 VSS 0.444691f
C9644 a_33812_n15304 VSS 0.442676f
C9645 a_33364_n15304 VSS 0.44117f
C9646 a_32916_n15304 VSS 0.480946f
C9647 a_27316_n14820 VSS 0.178831f
C9648 a_24116_n15216 VSS 0.012971f
C9649 a_25472_n14816 VSS 0.145471f
C9650 a_27852_n14990 VSS 0.814313f
C9651 a_27404_n14990 VSS 0.828568f
C9652 a_25160_n14816 VSS 0.380744f
C9653 a_25577_n14956 VSS 0.771187f
C9654 a_23912_n15216 VSS 0.335295f
C9655 a_23708_n15216 VSS 0.075356f
C9656 a_24220_n15260 VSS 0.280893f
C9657 a_23608_n15260 VSS 0.612054f
C9658 a_23360_n15233 VSS 1.87054f
C9659 a_22140_n15348 VSS 0.239647f
C9660 a_21692_n15348 VSS 0.295123f
C9661 a_22948_n14820 VSS 1.42665f
C9662 a_22052_n15304 VSS 0.462457f
C9663 a_21604_n15304 VSS 0.4881f
C9664 a_47924_n14116 VSS 0.474295f
C9665 a_47476_n14116 VSS 0.461553f
C9666 a_47028_n14116 VSS 0.45987f
C9667 a_46580_n14116 VSS 0.457171f
C9668 a_46132_n14116 VSS 0.45666f
C9669 a_45684_n14116 VSS 0.45666f
C9670 a_45236_n14116 VSS 0.45666f
C9671 a_44788_n14116 VSS 0.471552f
C9672 a_44340_n14116 VSS 0.457943f
C9673 a_43892_n14116 VSS 0.4579f
C9674 a_43444_n14116 VSS 0.458658f
C9675 a_42996_n14116 VSS 0.46122f
C9676 a_42548_n14116 VSS 0.463019f
C9677 a_42100_n14116 VSS 0.46578f
C9678 a_41652_n14116 VSS 0.499395f
C9679 a_41204_n14116 VSS 0.47766f
C9680 a_40532_n14116 VSS 0.474856f
C9681 a_40084_n14116 VSS 0.459483f
C9682 a_39636_n14116 VSS 0.45666f
C9683 a_39188_n14116 VSS 0.45666f
C9684 a_38740_n14116 VSS 0.45666f
C9685 a_38292_n14116 VSS 0.45666f
C9686 a_37844_n14116 VSS 0.45666f
C9687 a_37396_n14116 VSS 0.45666f
C9688 a_36948_n14116 VSS 0.471552f
C9689 a_36500_n14116 VSS 0.442251f
C9690 a_36052_n14116 VSS 0.443851f
C9691 a_35604_n14116 VSS 0.445739f
C9692 a_35156_n14116 VSS 0.446903f
C9693 a_34708_n14116 VSS 0.470374f
C9694 a_34260_n14116 VSS 0.446699f
C9695 a_33812_n14116 VSS 0.444684f
C9696 a_33364_n14116 VSS 0.455478f
C9697 a_48012_n14213 VSS 0.321039f
C9698 a_47564_n14213 VSS 0.290098f
C9699 a_47116_n14213 VSS 0.288045f
C9700 a_46668_n14213 VSS 0.28552f
C9701 a_46220_n14213 VSS 0.284099f
C9702 a_45772_n14213 VSS 0.284099f
C9703 a_45324_n14213 VSS 0.284099f
C9704 a_44876_n14213 VSS 0.285753f
C9705 a_44428_n14213 VSS 0.284269f
C9706 a_43980_n14213 VSS 0.284258f
C9707 a_43532_n14213 VSS 0.284258f
C9708 a_43084_n14213 VSS 0.287629f
C9709 a_42636_n14213 VSS 0.289343f
C9710 a_42188_n14213 VSS 0.290362f
C9711 a_41740_n14213 VSS 0.314383f
C9712 a_41292_n14213 VSS 0.298098f
C9713 a_40620_n14213 VSS 0.296372f
C9714 a_40172_n14213 VSS 0.292759f
C9715 a_39724_n14213 VSS 0.285905f
C9716 a_39276_n14213 VSS 0.285816f
C9717 a_38828_n14213 VSS 0.285815f
C9718 a_38380_n14213 VSS 0.285815f
C9719 a_37932_n14213 VSS 0.285815f
C9720 a_37484_n14213 VSS 0.285815f
C9721 a_37036_n14213 VSS 0.288747f
C9722 a_36588_n14213 VSS 0.283621f
C9723 a_36140_n14213 VSS 0.285724f
C9724 a_35692_n14213 VSS 0.287452f
C9725 a_35244_n14213 VSS 0.28974f
C9726 a_34796_n14213 VSS 0.325726f
C9727 a_34348_n14213 VSS 0.296215f
C9728 a_33900_n14213 VSS 0.290144f
C9729 a_33452_n14213 VSS 0.288574f
C9730 a_32413_n14564 VSS 0.768248f
C9731 a_31789_n14564 VSS 0.761795f
C9732 a_28752_n15348 VSS 1.80699f
C9733 a_31459_n14564 VSS 0.62655f
C9734 a_25636_n14520 VSS 0.183324f
C9735 a_29056_n14432 VSS 0.146547f
C9736 a_29161_n14476 VSS 0.772209f
C9737 a_28744_n14432 VSS 0.377456f
C9738 a_27700_n14116 VSS 0.020998f
C9739 a_27496_n14116 VSS 0.34666f
C9740 a_27292_n14116 VSS 0.076062f
C9741 a_27804_n14165 VSS 0.294505f
C9742 a_27192_n14286 VSS 0.597777f
C9743 a_26944_n14116 VSS 1.88836f
C9744 a_26532_n14437 VSS 1.40595f
C9745 a_24516_n14475 VSS 0.437044f
C9746 a_32412_n13648 VSS 0.012971f
C9747 a_47900_n13780 VSS 0.300977f
C9748 a_47452_n13780 VSS 0.294024f
C9749 a_47004_n13780 VSS 0.29129f
C9750 a_46556_n13780 VSS 0.287668f
C9751 a_46108_n13780 VSS 0.285997f
C9752 a_45660_n13780 VSS 0.285997f
C9753 a_45212_n13780 VSS 0.289177f
C9754 a_47812_n13736 VSS 0.483823f
C9755 a_47364_n13736 VSS 0.46949f
C9756 a_46916_n13736 VSS 0.46798f
C9757 a_46468_n13736 VSS 0.461248f
C9758 a_46020_n13736 VSS 0.461248f
C9759 a_45572_n13736 VSS 0.461248f
C9760 a_45124_n13736 VSS 0.473068f
C9761 a_44540_n13780 VSS 0.289463f
C9762 a_44092_n13780 VSS 0.287579f
C9763 a_43644_n13780 VSS 0.284099f
C9764 a_43196_n13780 VSS 0.287148f
C9765 a_42748_n13780 VSS 0.288687f
C9766 a_42300_n13780 VSS 0.28953f
C9767 a_41852_n13780 VSS 0.300321f
C9768 a_41404_n13780 VSS 0.308618f
C9769 a_40956_n13780 VSS 0.292892f
C9770 a_40508_n13780 VSS 0.289019f
C9771 a_40060_n13780 VSS 0.287384f
C9772 a_39612_n13780 VSS 0.284258f
C9773 a_39164_n13780 VSS 0.284258f
C9774 a_38716_n13780 VSS 0.284258f
C9775 a_38268_n13780 VSS 0.284258f
C9776 a_37820_n13780 VSS 0.284258f
C9777 a_37372_n13780 VSS 0.287991f
C9778 a_44452_n13736 VSS 0.470565f
C9779 a_44004_n13736 VSS 0.45666f
C9780 a_43556_n13736 VSS 0.45666f
C9781 a_43108_n13736 VSS 0.459647f
C9782 a_42660_n13736 VSS 0.461258f
C9783 a_42212_n13736 VSS 0.462696f
C9784 a_41764_n13736 VSS 0.485271f
C9785 a_41316_n13736 VSS 0.465969f
C9786 a_40868_n13736 VSS 0.477382f
C9787 a_40420_n13736 VSS 0.460519f
C9788 a_39972_n13736 VSS 0.458997f
C9789 a_39524_n13736 VSS 0.45666f
C9790 a_39076_n13736 VSS 0.45666f
C9791 a_38628_n13736 VSS 0.45666f
C9792 a_38180_n13736 VSS 0.45666f
C9793 a_37732_n13736 VSS 0.45666f
C9794 a_37284_n13736 VSS 0.471163f
C9795 a_36588_n13780 VSS 0.272289f
C9796 a_36140_n13780 VSS 0.289561f
C9797 a_35692_n13780 VSS 0.289861f
C9798 a_35244_n13780 VSS 0.292335f
C9799 a_34796_n13780 VSS 0.33077f
C9800 a_33280_n13248 VSS 0.076267f
C9801 a_36500_n13736 VSS 0.488036f
C9802 a_36052_n13736 VSS 0.479285f
C9803 a_35604_n13736 VSS 0.481308f
C9804 a_35156_n13736 VSS 0.482667f
C9805 a_34708_n13736 VSS 0.530158f
C9806 a_29479_n13735 VSS 0.028065f
C9807 a_31960_n13648 VSS 0.282998f
C9808 a_31455_n13648 VSS 0.145471f
C9809 a_32152_n13692 VSS 0.33544f
C9810 a_31559_n13692 VSS 1.87864f
C9811 a_31664_n13292 VSS 1.44889f
C9812 a_30903_n13780 VSS 0.388656f
C9813 a_27820_n16432 VSS 0.812861f
C9814 a_30555_n13780 VSS 0.75771f
C9815 a_30159_n13296 VSS 0.560529f
C9816 a_22772_n13648 VSS 0.012971f
C9817 a_24128_n13248 VSS 0.145471f
C9818 a_27526_n13714 VSS 0.667711f
C9819 a_27302_n13160 VSS 0.728255f
C9820 a_26470_n13736 VSS 0.934072f
C9821 a_26266_n13736 VSS 0.742882f
C9822 a_25642_n13736 VSS 0.729211f
C9823 a_25237_n13735 VSS 0.722244f
C9824 a_23816_n13248 VSS 0.368907f
C9825 a_24233_n13388 VSS 0.77136f
C9826 a_22568_n13648 VSS 0.335295f
C9827 a_22364_n13648 VSS 0.075356f
C9828 a_22876_n13692 VSS 0.288657f
C9829 a_22016_n13665 VSS 1.8736f
C9830 a_21604_n13252 VSS 1.42418f
C9831 a_47924_n12548 VSS 0.474295f
C9832 a_47476_n12548 VSS 0.461553f
C9833 a_47028_n12548 VSS 0.45987f
C9834 a_46580_n12548 VSS 0.457171f
C9835 a_46132_n12548 VSS 0.45666f
C9836 a_45684_n12548 VSS 0.45666f
C9837 a_45236_n12548 VSS 0.45666f
C9838 a_44788_n12548 VSS 0.471552f
C9839 a_44340_n12548 VSS 0.457943f
C9840 a_43892_n12548 VSS 0.4579f
C9841 a_43444_n12548 VSS 0.458658f
C9842 a_42996_n12548 VSS 0.46122f
C9843 a_42548_n12548 VSS 0.463019f
C9844 a_42100_n12548 VSS 0.46578f
C9845 a_41652_n12548 VSS 0.499395f
C9846 a_41204_n12548 VSS 0.482015f
C9847 a_40308_n12548 VSS 0.476821f
C9848 a_39860_n12548 VSS 0.467616f
C9849 a_39412_n12548 VSS 0.466435f
C9850 a_38964_n12548 VSS 0.462598f
C9851 a_38516_n12548 VSS 0.462598f
C9852 a_38068_n12548 VSS 0.462598f
C9853 a_37620_n12548 VSS 0.462598f
C9854 a_37172_n12548 VSS 0.457242f
C9855 a_36724_n12548 VSS 0.469961f
C9856 a_36276_n12548 VSS 0.47378f
C9857 a_35828_n12548 VSS 0.475941f
C9858 a_35380_n12548 VSS 0.47834f
C9859 a_34932_n12548 VSS 0.500343f
C9860 a_34484_n12548 VSS 0.47638f
C9861 a_34036_n12548 VSS 0.476399f
C9862 a_48012_n12645 VSS 0.321039f
C9863 a_47564_n12645 VSS 0.290098f
C9864 a_47116_n12645 VSS 0.288045f
C9865 a_46668_n12645 VSS 0.28552f
C9866 a_46220_n12645 VSS 0.284099f
C9867 a_45772_n12645 VSS 0.284099f
C9868 a_45324_n12645 VSS 0.284099f
C9869 a_44876_n12645 VSS 0.285753f
C9870 a_44428_n12645 VSS 0.284269f
C9871 a_43980_n12645 VSS 0.284258f
C9872 a_43532_n12645 VSS 0.284258f
C9873 a_43084_n12645 VSS 0.287629f
C9874 a_42636_n12645 VSS 0.289343f
C9875 a_42188_n12645 VSS 0.290362f
C9876 a_41740_n12645 VSS 0.314383f
C9877 a_41292_n12645 VSS 0.298511f
C9878 a_40396_n12645 VSS 0.275298f
C9879 a_39948_n12645 VSS 0.292609f
C9880 a_39500_n12645 VSS 0.289367f
C9881 a_39052_n12645 VSS 0.288933f
C9882 a_38604_n12645 VSS 0.287628f
C9883 a_38156_n12645 VSS 0.287628f
C9884 a_37708_n12645 VSS 0.287628f
C9885 a_37260_n12645 VSS 0.286904f
C9886 a_36812_n12645 VSS 0.284653f
C9887 a_36364_n12645 VSS 0.287077f
C9888 a_35916_n12645 VSS 0.289278f
C9889 a_35468_n12645 VSS 0.29149f
C9890 a_35020_n12645 VSS 0.295434f
C9891 a_34572_n12645 VSS 0.299006f
C9892 a_34124_n12645 VSS 0.284985f
C9893 a_33488_n12996 VSS 0.365077f
C9894 a_32413_n12996 VSS 0.746281f
C9895 a_31789_n12996 VSS 0.73555f
C9896 a_29360_n12864 VSS 0.075356f
C9897 a_30340_n12548 VSS 0.480039f
C9898 a_31459_n12996 VSS 0.616954f
C9899 a_30428_n12645 VSS 0.240559f
C9900 a_28492_n12548 VSS 0.014625f
C9901 a_28040_n12493 VSS 0.311202f
C9902 a_27535_n12493 VSS 0.147013f
C9903 a_28232_n12606 VSS 0.345965f
C9904 a_27639_n12537 VSS 1.90773f
C9905 a_25132_n16432 VSS 0.744047f
C9906 a_25559_n12548 VSS 0.026839f
C9907 a_21892_n12952 VSS 0.15997f
C9908 a_27744_n12908 VSS 1.46524f
C9909 a_26983_n12728 VSS 0.381013f
C9910 a_26635_n12996 VSS 0.753745f
C9911 a_26239_n12996 VSS 0.732f
C9912 a_25831_n12996 VSS 1.31572f
C9913 a_24573_n12996 VSS 0.761852f
C9914 a_23949_n12996 VSS 0.732104f
C9915 a_22264_n13692 VSS 0.616218f
C9916 a_21872_n12530 VSS 0.693301f
C9917 a_23619_n12996 VSS 0.616146f
C9918 a_21772_n12996 VSS 1.70852f
C9919 a_47900_n12212 VSS 0.300977f
C9920 a_47452_n12212 VSS 0.294024f
C9921 a_47004_n12212 VSS 0.29129f
C9922 a_46556_n12212 VSS 0.287668f
C9923 a_46108_n12212 VSS 0.285997f
C9924 a_45660_n12212 VSS 0.285997f
C9925 a_45212_n12212 VSS 0.289177f
C9926 a_47812_n12168 VSS 0.483823f
C9927 a_47364_n12168 VSS 0.46949f
C9928 a_46916_n12168 VSS 0.46798f
C9929 a_46468_n12168 VSS 0.461248f
C9930 a_46020_n12168 VSS 0.461248f
C9931 a_45572_n12168 VSS 0.461248f
C9932 a_45124_n12168 VSS 0.473068f
C9933 a_44540_n12212 VSS 0.289463f
C9934 a_44092_n12212 VSS 0.287579f
C9935 a_43644_n12212 VSS 0.284099f
C9936 a_43196_n12212 VSS 0.287148f
C9937 a_42748_n12212 VSS 0.288687f
C9938 a_42300_n12212 VSS 0.28953f
C9939 a_41852_n12212 VSS 0.300321f
C9940 a_41404_n12212 VSS 0.308618f
C9941 a_40956_n12212 VSS 0.292892f
C9942 a_40508_n12212 VSS 0.28885f
C9943 a_40060_n12212 VSS 0.287225f
C9944 a_39612_n12212 VSS 0.284099f
C9945 a_39164_n12212 VSS 0.284099f
C9946 a_38716_n12212 VSS 0.284099f
C9947 a_38268_n12212 VSS 0.284099f
C9948 a_37820_n12212 VSS 0.284099f
C9949 a_37372_n12212 VSS 0.2876f
C9950 a_44452_n12168 VSS 0.470565f
C9951 a_44004_n12168 VSS 0.45666f
C9952 a_43556_n12168 VSS 0.45666f
C9953 a_43108_n12168 VSS 0.459647f
C9954 a_42660_n12168 VSS 0.461258f
C9955 a_42212_n12168 VSS 0.462696f
C9956 a_41764_n12168 VSS 0.485271f
C9957 a_41316_n12168 VSS 0.465969f
C9958 a_40868_n12168 VSS 0.477382f
C9959 a_40420_n12168 VSS 0.461791f
C9960 a_39972_n12168 VSS 0.460269f
C9961 a_39524_n12168 VSS 0.457889f
C9962 a_39076_n12168 VSS 0.457889f
C9963 a_38628_n12168 VSS 0.457889f
C9964 a_38180_n12168 VSS 0.457889f
C9965 a_37732_n12168 VSS 0.457889f
C9966 a_37284_n12168 VSS 0.469849f
C9967 a_36700_n12212 VSS 0.289363f
C9968 a_36252_n12212 VSS 0.2883f
C9969 a_35804_n12212 VSS 0.290851f
C9970 a_35356_n12212 VSS 0.29392f
C9971 a_30599_n12167 VSS 0.026799f
C9972 a_31760_n12168 VSS 0.747658f
C9973 a_30787_n12167 VSS 0.542553f
C9974 a_36612_n12168 VSS 0.466184f
C9975 a_36164_n12168 VSS 0.476489f
C9976 a_35716_n12168 VSS 0.479839f
C9977 a_35268_n12168 VSS 0.492582f
C9978 a_33910_n12146 VSS 0.66738f
C9979 a_33686_n11592 VSS 0.763756f
C9980 a_32854_n12168 VSS 0.943593f
C9981 a_32650_n12168 VSS 0.759811f
C9982 a_32026_n12168 VSS 0.727934f
C9983 a_31279_n11728 VSS 0.41599f
C9984 a_29540_n11728 VSS 0.980011f
C9985 a_28009_n12168 VSS 0.612767f
C9986 a_25880_n11708 VSS 0.410111f
C9987 a_23108_n12080 VSS 0.012971f
C9988 a_24464_n11680 VSS 0.145471f
C9989 a_27279_n12146 VSS 0.646359f
C9990 a_27055_n12168 VSS 0.763947f
C9991 a_26431_n12168 VSS 0.730957f
C9992 a_26563_n12212 VSS 0.811729f
C9993 a_24152_n11680 VSS 0.380215f
C9994 a_24569_n11820 VSS 0.771138f
C9995 a_22904_n12080 VSS 0.335295f
C9996 a_22700_n12080 VSS 0.075356f
C9997 a_23212_n12124 VSS 0.286776f
C9998 a_22600_n12124 VSS 0.926517f
C9999 a_22352_n12097 VSS 1.86892f
C10000 a_21940_n11684 VSS 1.41883f
C10001 a_47924_n10980 VSS 0.474295f
C10002 a_47476_n10980 VSS 0.461553f
C10003 a_47028_n10980 VSS 0.45987f
C10004 a_46580_n10980 VSS 0.457171f
C10005 a_46132_n10980 VSS 0.45666f
C10006 a_45684_n10980 VSS 0.45666f
C10007 a_45236_n10980 VSS 0.45666f
C10008 a_44788_n10980 VSS 0.471552f
C10009 a_44340_n10980 VSS 0.457943f
C10010 a_43892_n10980 VSS 0.4579f
C10011 a_43444_n10980 VSS 0.458658f
C10012 a_42996_n10980 VSS 0.46122f
C10013 a_42548_n10980 VSS 0.463019f
C10014 a_42100_n10980 VSS 0.46578f
C10015 a_41652_n10980 VSS 0.499395f
C10016 a_41204_n10980 VSS 0.47766f
C10017 a_40532_n10980 VSS 0.473316f
C10018 a_40084_n10980 VSS 0.468056f
C10019 a_39636_n10980 VSS 0.45604f
C10020 a_39188_n10980 VSS 0.45604f
C10021 a_38740_n10980 VSS 0.456039f
C10022 a_38292_n10980 VSS 0.456039f
C10023 a_37844_n10980 VSS 0.456039f
C10024 a_37396_n10980 VSS 0.456039f
C10025 a_36948_n10980 VSS 0.471991f
C10026 a_33364_n11384 VSS 0.200437f
C10027 a_36500_n10980 VSS 0.483406f
C10028 a_28300_n15348 VSS 1.8147f
C10029 a_32158_n12212 VSS 0.865894f
C10030 a_48012_n11077 VSS 0.321039f
C10031 a_47564_n11077 VSS 0.290098f
C10032 a_47116_n11077 VSS 0.288045f
C10033 a_46668_n11077 VSS 0.28552f
C10034 a_46220_n11077 VSS 0.284099f
C10035 a_45772_n11077 VSS 0.284099f
C10036 a_45324_n11077 VSS 0.284099f
C10037 a_44876_n11077 VSS 0.285753f
C10038 a_44428_n11077 VSS 0.284269f
C10039 a_43980_n11077 VSS 0.284258f
C10040 a_43532_n11077 VSS 0.284258f
C10041 a_43084_n11077 VSS 0.287629f
C10042 a_42636_n11077 VSS 0.289343f
C10043 a_42188_n11077 VSS 0.290362f
C10044 a_41740_n11077 VSS 0.314383f
C10045 a_41292_n11077 VSS 0.298098f
C10046 a_40620_n11077 VSS 0.294453f
C10047 a_40172_n11077 VSS 0.29104f
C10048 a_39724_n11077 VSS 0.286509f
C10049 a_39276_n11077 VSS 0.28294f
C10050 a_38828_n11077 VSS 0.28294f
C10051 a_38380_n11077 VSS 0.28294f
C10052 a_37932_n11077 VSS 0.28294f
C10053 a_37484_n11077 VSS 0.28294f
C10054 a_37036_n11077 VSS 0.284593f
C10055 a_36588_n11077 VSS 0.28599f
C10056 a_34350_n10980 VSS 0.732437f
C10057 a_35064_n11383 VSS 0.442524f
C10058 a_31856_n11296 VSS 0.145471f
C10059 a_31961_n11340 VSS 0.769349f
C10060 a_31544_n11296 VSS 0.373304f
C10061 a_30500_n10980 VSS 0.012971f
C10062 a_30296_n10980 VSS 0.335295f
C10063 a_30092_n10980 VSS 0.075356f
C10064 a_30604_n11029 VSS 0.285207f
C10065 a_29744_n10980 VSS 1.873f
C10066 a_28121_n10980 VSS 1.28608f
C10067 a_29332_n11301 VSS 1.43413f
C10068 a_27391_n11384 VSS 0.667143f
C10069 a_27167_n10808 VSS 0.758019f
C10070 a_24684_n16432 VSS 0.758743f
C10071 a_25559_n10980 VSS 0.026878f
C10072 a_26543_n11384 VSS 0.733748f
C10073 a_26547_n12951 VSS 0.769701f
C10074 a_24964_n14116 VSS 2.03276f
C10075 a_24760_n11383 VSS 0.456773f
C10076 a_23564_n11428 VSS 1.65805f
C10077 a_47900_n10644 VSS 0.300977f
C10078 a_47452_n10644 VSS 0.294024f
C10079 a_47004_n10644 VSS 0.29129f
C10080 a_46556_n10644 VSS 0.287668f
C10081 a_46108_n10644 VSS 0.285997f
C10082 a_45660_n10644 VSS 0.285997f
C10083 a_45212_n10644 VSS 0.289177f
C10084 a_47812_n10600 VSS 0.483823f
C10085 a_47364_n10600 VSS 0.46949f
C10086 a_46916_n10600 VSS 0.46798f
C10087 a_46468_n10600 VSS 0.461248f
C10088 a_46020_n10600 VSS 0.461248f
C10089 a_45572_n10600 VSS 0.461248f
C10090 a_45124_n10600 VSS 0.473068f
C10091 a_44540_n10644 VSS 0.289463f
C10092 a_44092_n10644 VSS 0.287579f
C10093 a_43644_n10644 VSS 0.284099f
C10094 a_43196_n10644 VSS 0.287148f
C10095 a_42748_n10644 VSS 0.288687f
C10096 a_42300_n10644 VSS 0.28953f
C10097 a_41852_n10644 VSS 0.300321f
C10098 a_41404_n10644 VSS 0.308618f
C10099 a_40956_n10644 VSS 0.292892f
C10100 a_40508_n10644 VSS 0.289017f
C10101 a_40060_n10644 VSS 0.287391f
C10102 a_39612_n10644 VSS 0.284256f
C10103 a_39164_n10644 VSS 0.284256f
C10104 a_38716_n10644 VSS 0.284256f
C10105 a_38268_n10644 VSS 0.284256f
C10106 a_37820_n10644 VSS 0.284256f
C10107 a_37372_n10644 VSS 0.288286f
C10108 a_44452_n10600 VSS 0.470565f
C10109 a_44004_n10600 VSS 0.45666f
C10110 a_43556_n10600 VSS 0.45666f
C10111 a_43108_n10600 VSS 0.459647f
C10112 a_42660_n10600 VSS 0.461258f
C10113 a_42212_n10600 VSS 0.462696f
C10114 a_41764_n10600 VSS 0.485271f
C10115 a_41316_n10600 VSS 0.465969f
C10116 a_40868_n10600 VSS 0.477382f
C10117 a_40420_n10600 VSS 0.461791f
C10118 a_39972_n10600 VSS 0.460269f
C10119 a_39524_n10600 VSS 0.457889f
C10120 a_39076_n10600 VSS 0.457889f
C10121 a_38628_n10600 VSS 0.457889f
C10122 a_38180_n10600 VSS 0.457889f
C10123 a_37732_n10600 VSS 0.457889f
C10124 a_37284_n10600 VSS 0.475005f
C10125 a_33900_n11428 VSS 0.799837f
C10126 a_34652_n11391 VSS 1.16093f
C10127 a_32628_n10512 VSS 0.013111f
C10128 a_33984_n10112 VSS 0.146478f
C10129 a_30871_n11728 VSS 1.45362f
C10130 a_35392_n10172 VSS 0.354875f
C10131 a_33672_n10112 VSS 0.387176f
C10132 a_34089_n10252 VSS 0.789145f
C10133 a_32424_n10512 VSS 0.336354f
C10134 a_32220_n10512 VSS 0.075356f
C10135 a_32732_n10556 VSS 0.291888f
C10136 a_31872_n10529 VSS 1.87025f
C10137 a_30808_n10116 VSS 0.666918f
C10138 a_28247_n10599 VSS 0.036737f
C10139 a_31460_n10116 VSS 1.40215f
C10140 a_30136_n10600 VSS 0.715356f
C10141 a_29444_n10116 VSS 0.377641f
C10142 a_28435_n10599 VSS 0.452847f
C10143 a_28927_n10160 VSS 1.73304f
C10144 a_28437_n13705 VSS 0.604099f
C10145 a_26239_n11428 VSS 0.476335f
C10146 a_25500_n10644 VSS 0.240066f
C10147 a_22772_n10512 VSS 0.012971f
C10148 a_24128_n10112 VSS 0.145471f
C10149 a_27485_n10068 VSS 0.772473f
C10150 a_26861_n10135 VSS 0.747185f
C10151 a_26531_n10207 VSS 0.630485f
C10152 a_25412_n10600 VSS 0.483018f
C10153 a_23816_n10112 VSS 0.368329f
C10154 a_24233_n10252 VSS 0.768713f
C10155 a_22568_n10512 VSS 0.335295f
C10156 a_22364_n10512 VSS 0.075356f
C10157 a_22876_n10556 VSS 0.288657f
C10158 a_22016_n10529 VSS 1.8736f
C10159 a_21604_n10116 VSS 1.42231f
C10160 a_47924_n9412 VSS 0.474295f
C10161 a_47476_n9412 VSS 0.461553f
C10162 a_47028_n9412 VSS 0.45987f
C10163 a_46580_n9412 VSS 0.457171f
C10164 a_46132_n9412 VSS 0.45666f
C10165 a_45684_n9412 VSS 0.45666f
C10166 a_45236_n9412 VSS 0.45666f
C10167 a_44788_n9412 VSS 0.471552f
C10168 a_44340_n9412 VSS 0.457943f
C10169 a_43892_n9412 VSS 0.4579f
C10170 a_43444_n9412 VSS 0.458658f
C10171 a_42996_n9412 VSS 0.46122f
C10172 a_42548_n9412 VSS 0.463019f
C10173 a_42100_n9412 VSS 0.46578f
C10174 a_41652_n9412 VSS 0.499395f
C10175 a_41204_n9412 VSS 0.47766f
C10176 a_40532_n9412 VSS 0.471965f
C10177 a_40084_n9412 VSS 0.466668f
C10178 a_39636_n9412 VSS 0.454653f
C10179 a_39188_n9412 VSS 0.454653f
C10180 a_38740_n9412 VSS 0.454653f
C10181 a_38292_n9412 VSS 0.454653f
C10182 a_37844_n9412 VSS 0.454653f
C10183 a_37396_n9412 VSS 0.454653f
C10184 a_36948_n9412 VSS 0.469545f
C10185 a_36500_n9412 VSS 0.494161f
C10186 a_25020_n11383 VSS 1.22928f
C10187 a_28335_n10644 VSS 0.821665f
C10188 a_48012_n9509 VSS 0.321039f
C10189 a_47564_n9509 VSS 0.290098f
C10190 a_47116_n9509 VSS 0.288045f
C10191 a_46668_n9509 VSS 0.28552f
C10192 a_46220_n9509 VSS 0.284099f
C10193 a_45772_n9509 VSS 0.284099f
C10194 a_45324_n9509 VSS 0.284099f
C10195 a_44876_n9509 VSS 0.285753f
C10196 a_44428_n9509 VSS 0.284269f
C10197 a_43980_n9509 VSS 0.284258f
C10198 a_43532_n9509 VSS 0.284258f
C10199 a_43084_n9509 VSS 0.287629f
C10200 a_42636_n9509 VSS 0.289343f
C10201 a_42188_n9509 VSS 0.290362f
C10202 a_41740_n9509 VSS 0.314383f
C10203 a_41292_n9509 VSS 0.298098f
C10204 a_40620_n9509 VSS 0.296083f
C10205 a_40172_n9509 VSS 0.292756f
C10206 a_39724_n9509 VSS 0.288226f
C10207 a_39276_n9509 VSS 0.284653f
C10208 a_38828_n9509 VSS 0.284653f
C10209 a_38380_n9509 VSS 0.284653f
C10210 a_37932_n9509 VSS 0.284653f
C10211 a_37484_n9509 VSS 0.284653f
C10212 a_37036_n9509 VSS 0.287587f
C10213 a_36588_n9509 VSS 0.289188f
C10214 a_34392_n9815 VSS 0.463975f
C10215 a_33494_n9860 VSS 0.694066f
C10216 a_32581_n9860 VSS 0.751398f
C10217 a_32189_n9860 VSS 0.731055f
C10218 a_31565_n9860 VSS 0.75622f
C10219 a_29992_n11150 VSS 0.530574f
C10220 a_25724_n14564 VSS 1.31249f
C10221 a_28644_n9815 VSS 0.710077f
C10222 a_22220_n12996 VSS 1.17528f
C10223 a_31235_n9860 VSS 0.633112f
C10224 a_30472_n9815 VSS 0.417675f
C10225 a_28624_n9394 VSS 0.562006f
C10226 a_29800_n9815 VSS 0.405125f
C10227 a_27281_n16854 VSS 1.08199f
C10228 a_27526_n9816 VSS 0.692245f
C10229 a_27302_n9816 VSS 0.729716f
C10230 a_21892_n9816 VSS 0.1641f
C10231 a_26470_n9322 VSS 0.938441f
C10232 a_26266_n9240 VSS 0.74647f
C10233 a_25642_n9816 VSS 0.776211f
C10234 a_25237_n10599 VSS 0.807507f
C10235 a_24965_n9860 VSS 0.856529f
C10236 a_24573_n9860 VSS 0.762883f
C10237 a_23949_n9860 VSS 0.732356f
C10238 a_22264_n10556 VSS 0.608542f
C10239 a_23619_n9860 VSS 0.616146f
C10240 a_21772_n9860 VSS 1.09751f
C10241 a_47900_n9076 VSS 0.300977f
C10242 a_47452_n9076 VSS 0.294024f
C10243 a_47004_n9076 VSS 0.29129f
C10244 a_46556_n9076 VSS 0.287668f
C10245 a_46108_n9076 VSS 0.285997f
C10246 a_45660_n9076 VSS 0.285997f
C10247 a_45212_n9076 VSS 0.289177f
C10248 a_47812_n9032 VSS 0.483823f
C10249 a_47364_n9032 VSS 0.46949f
C10250 a_46916_n9032 VSS 0.46798f
C10251 a_46468_n9032 VSS 0.461248f
C10252 a_46020_n9032 VSS 0.461248f
C10253 a_45572_n9032 VSS 0.461248f
C10254 a_45124_n9032 VSS 0.473068f
C10255 a_44540_n9076 VSS 0.289463f
C10256 a_44092_n9076 VSS 0.287579f
C10257 a_43644_n9076 VSS 0.284099f
C10258 a_43196_n9076 VSS 0.287148f
C10259 a_42748_n9076 VSS 0.288687f
C10260 a_42300_n9076 VSS 0.28953f
C10261 a_41852_n9076 VSS 0.300321f
C10262 a_41404_n9076 VSS 0.308618f
C10263 a_40956_n9076 VSS 0.292892f
C10264 a_40508_n9076 VSS 0.289017f
C10265 a_40060_n9076 VSS 0.287391f
C10266 a_39612_n9076 VSS 0.284256f
C10267 a_39164_n9076 VSS 0.284256f
C10268 a_38716_n9076 VSS 0.284256f
C10269 a_38268_n9076 VSS 0.284256f
C10270 a_37820_n9076 VSS 0.284256f
C10271 a_37372_n9076 VSS 0.288286f
C10272 a_44452_n9032 VSS 0.470565f
C10273 a_44004_n9032 VSS 0.45666f
C10274 a_43556_n9032 VSS 0.45666f
C10275 a_43108_n9032 VSS 0.459647f
C10276 a_42660_n9032 VSS 0.461258f
C10277 a_42212_n9032 VSS 0.462696f
C10278 a_41764_n9032 VSS 0.485271f
C10279 a_41316_n9032 VSS 0.465969f
C10280 a_40868_n9032 VSS 0.477382f
C10281 a_40420_n9032 VSS 0.460519f
C10282 a_39972_n9032 VSS 0.458997f
C10283 a_39524_n9032 VSS 0.45666f
C10284 a_39076_n9032 VSS 0.45666f
C10285 a_38628_n9032 VSS 0.45666f
C10286 a_38180_n9032 VSS 0.45666f
C10287 a_37732_n9032 VSS 0.45666f
C10288 a_37284_n9032 VSS 0.473776f
C10289 a_25831_n11428 VSS 1.33143f
C10290 a_34092_n9076 VSS 0.662088f
C10291 a_33832_n8572 VSS 0.450032f
C10292 a_28225_n9031 VSS 0.040346f
C10293 a_32767_n9010 VSS 0.634294f
C10294 a_32543_n9032 VSS 0.765641f
C10295 a_31919_n9032 VSS 0.742408f
C10296 a_30900_n9032 VSS 0.712949f
C10297 a_28617_n8548 VSS 0.493158f
C10298 a_25573_n12167 VSS 1.99485f
C10299 a_25860_n9032 VSS 0.752115f
C10300 a_25412_n8501 VSS 0.414925f
C10301 a_22772_n8944 VSS 0.012971f
C10302 a_24128_n8544 VSS 0.145471f
C10303 a_21872_n9394 VSS 0.782546f
C10304 a_27485_n8500 VSS 0.769614f
C10305 a_26861_n8567 VSS 0.759312f
C10306 a_26531_n8639 VSS 0.632421f
C10307 a_23816_n8544 VSS 0.366362f
C10308 a_24233_n8684 VSS 0.769723f
C10309 a_22568_n8944 VSS 0.335295f
C10310 a_22364_n8944 VSS 0.075356f
C10311 a_22876_n8988 VSS 0.280882f
C10312 a_22264_n8988 VSS 0.726892f
C10313 a_22016_n8961 VSS 1.86843f
C10314 a_21604_n8548 VSS 1.43225f
C10315 a_47924_n7844 VSS 0.474295f
C10316 a_47476_n7844 VSS 0.461553f
C10317 a_47028_n7844 VSS 0.45987f
C10318 a_46580_n7844 VSS 0.457171f
C10319 a_46132_n7844 VSS 0.45666f
C10320 a_45684_n7844 VSS 0.45666f
C10321 a_45236_n7844 VSS 0.45666f
C10322 a_44788_n7844 VSS 0.471552f
C10323 a_44340_n7844 VSS 0.457943f
C10324 a_43892_n7844 VSS 0.4579f
C10325 a_43444_n7844 VSS 0.458658f
C10326 a_42996_n7844 VSS 0.46122f
C10327 a_42548_n7844 VSS 0.463019f
C10328 a_42100_n7844 VSS 0.46578f
C10329 a_41652_n7844 VSS 0.499395f
C10330 a_41204_n7844 VSS 0.482015f
C10331 a_40308_n7844 VSS 0.473931f
C10332 a_39860_n7844 VSS 0.467616f
C10333 a_39412_n7844 VSS 0.457242f
C10334 a_38964_n7844 VSS 0.457242f
C10335 a_38516_n7844 VSS 0.457242f
C10336 a_38068_n7844 VSS 0.457242f
C10337 a_37620_n7844 VSS 0.457242f
C10338 a_37172_n7844 VSS 0.457242f
C10339 a_36724_n7844 VSS 0.46996f
C10340 a_36276_n7844 VSS 0.488274f
C10341 a_29532_n10311 VSS 1.90058f
C10342 a_48012_n7941 VSS 0.321039f
C10343 a_47564_n7941 VSS 0.290098f
C10344 a_47116_n7941 VSS 0.288045f
C10345 a_46668_n7941 VSS 0.28552f
C10346 a_46220_n7941 VSS 0.284099f
C10347 a_45772_n7941 VSS 0.284099f
C10348 a_45324_n7941 VSS 0.284099f
C10349 a_44876_n7941 VSS 0.285753f
C10350 a_44428_n7941 VSS 0.284269f
C10351 a_43980_n7941 VSS 0.284258f
C10352 a_43532_n7941 VSS 0.284258f
C10353 a_43084_n7941 VSS 0.287629f
C10354 a_42636_n7941 VSS 0.289343f
C10355 a_42188_n7941 VSS 0.290362f
C10356 a_41740_n7941 VSS 0.314383f
C10357 a_41292_n7941 VSS 0.298511f
C10358 a_40396_n7941 VSS 0.273378f
C10359 a_39948_n7941 VSS 0.290109f
C10360 a_39500_n7941 VSS 0.286579f
C10361 a_39052_n7941 VSS 0.284729f
C10362 a_38604_n7941 VSS 0.283687f
C10363 a_38156_n7941 VSS 0.283579f
C10364 a_37708_n7941 VSS 0.283579f
C10365 a_37260_n7941 VSS 0.283579f
C10366 a_36812_n7941 VSS 0.285307f
C10367 a_36364_n7941 VSS 0.288118f
C10368 a_31965_n8292 VSS 0.731577f
C10369 a_31341_n8292 VSS 0.752265f
C10370 a_30676_n7844 VSS 0.784581f
C10371 a_28972_n8247 VSS 0.710008f
C10372 a_31011_n8292 VSS 0.618285f
C10373 a_30228_n8203 VSS 0.430133f
C10374 a_28764_n8247 VSS 0.585525f
C10375 a_27597_n8292 VSS 0.783545f
C10376 a_26973_n8292 VSS 0.759117f
C10377 a_26643_n8292 VSS 0.634157f
C10378 a_24752_n8292 VSS 0.373986f
C10379 a_23564_n8292 VSS 1.62599f
C10380 a_33308_n7376 VSS 0.01439f
C10381 a_47900_n7508 VSS 0.300977f
C10382 a_47452_n7508 VSS 0.294024f
C10383 a_47004_n7508 VSS 0.29129f
C10384 a_46556_n7508 VSS 0.287668f
C10385 a_46108_n7508 VSS 0.285997f
C10386 a_45660_n7508 VSS 0.285997f
C10387 a_45212_n7508 VSS 0.289177f
C10388 a_47812_n7464 VSS 0.483823f
C10389 a_47364_n7464 VSS 0.46949f
C10390 a_46916_n7464 VSS 0.46798f
C10391 a_46468_n7464 VSS 0.461248f
C10392 a_46020_n7464 VSS 0.461248f
C10393 a_45572_n7464 VSS 0.461248f
C10394 a_45124_n7464 VSS 0.473068f
C10395 a_44540_n7508 VSS 0.289463f
C10396 a_44092_n7508 VSS 0.287579f
C10397 a_43644_n7508 VSS 0.284099f
C10398 a_43196_n7508 VSS 0.287148f
C10399 a_42748_n7508 VSS 0.288687f
C10400 a_42300_n7508 VSS 0.28953f
C10401 a_41852_n7508 VSS 0.300321f
C10402 a_41404_n7508 VSS 0.308618f
C10403 a_40956_n7508 VSS 0.292892f
C10404 a_40508_n7508 VSS 0.28885f
C10405 a_40060_n7508 VSS 0.287225f
C10406 a_39612_n7508 VSS 0.284099f
C10407 a_39164_n7508 VSS 0.284099f
C10408 a_38716_n7508 VSS 0.284099f
C10409 a_38268_n7508 VSS 0.284099f
C10410 a_37820_n7508 VSS 0.284099f
C10411 a_37372_n7508 VSS 0.289057f
C10412 a_44452_n7464 VSS 0.471915f
C10413 a_44004_n7464 VSS 0.45695f
C10414 a_43556_n7464 VSS 0.45695f
C10415 a_43108_n7464 VSS 0.459937f
C10416 a_42660_n7464 VSS 0.461547f
C10417 a_42212_n7464 VSS 0.462985f
C10418 a_41764_n7464 VSS 0.48556f
C10419 a_41316_n7464 VSS 0.466249f
C10420 a_40868_n7464 VSS 0.478767f
C10421 a_40420_n7464 VSS 0.460808f
C10422 a_39972_n7464 VSS 0.459286f
C10423 a_39524_n7464 VSS 0.457289f
C10424 a_39076_n7464 VSS 0.471858f
C10425 a_38628_n7464 VSS 0.469369f
C10426 a_38180_n7464 VSS 0.464677f
C10427 a_37732_n7464 VSS 0.464677f
C10428 a_37284_n7464 VSS 0.482553f
C10429 a_34176_n6976 VSS 0.0771f
C10430 a_33497_n9032 VSS 0.552395f
C10431 a_32856_n7376 VSS 0.287446f
C10432 a_32351_n7376 VSS 0.145471f
C10433 a_33048_n7420 VSS 0.338317f
C10434 a_32455_n7420 VSS 1.88378f
C10435 a_32560_n7020 VSS 1.43751f
C10436 a_31799_n7508 VSS 0.370437f
C10437 a_31451_n7508 VSS 0.764077f
C10438 a_30036_n7464 VSS 1.0109f
C10439 a_30396_n7508 VSS 0.346318f
C10440 a_29476_n6980 VSS 0.458285f
C10441 a_23220_n7376 VSS 0.012971f
C10442 a_24576_n6976 VSS 0.145471f
C10443 a_26943_n7442 VSS 0.635074f
C10444 a_26719_n7464 VSS 0.762978f
C10445 a_26095_n7464 VSS 0.74528f
C10446 a_25685_n7463 VSS 0.714967f
C10447 a_24264_n6976 VSS 0.388135f
C10448 a_24681_n7116 VSS 0.765702f
C10449 a_23016_n7376 VSS 0.335295f
C10450 a_22812_n7376 VSS 0.075356f
C10451 a_23324_n7420 VSS 0.288403f
C10452 a_22712_n7420 VSS 0.534032f
C10453 a_22464_n7393 VSS 1.87233f
C10454 a_22052_n6980 VSS 1.41183f
C10455 a_47924_n6276 VSS 0.474295f
C10456 a_47476_n6276 VSS 0.461553f
C10457 a_47028_n6276 VSS 0.45987f
C10458 a_46580_n6276 VSS 0.457171f
C10459 a_46132_n6276 VSS 0.45666f
C10460 a_45684_n6276 VSS 0.45666f
C10461 a_45236_n6276 VSS 0.45666f
C10462 a_44788_n6276 VSS 0.471552f
C10463 a_44340_n6276 VSS 0.457943f
C10464 a_43892_n6276 VSS 0.4579f
C10465 a_43444_n6276 VSS 0.458658f
C10466 a_42996_n6276 VSS 0.46122f
C10467 a_42548_n6276 VSS 0.463019f
C10468 a_42100_n6276 VSS 0.464966f
C10469 a_41652_n6276 VSS 0.496709f
C10470 a_41204_n6276 VSS 0.481146f
C10471 a_40308_n6276 VSS 0.474995f
C10472 a_39860_n6276 VSS 0.466013f
C10473 a_39412_n6276 VSS 0.487547f
C10474 a_31936_n6592 VSS 0.075356f
C10475 a_48012_n6373 VSS 0.321039f
C10476 a_47564_n6373 VSS 0.290098f
C10477 a_47116_n6373 VSS 0.288045f
C10478 a_46668_n6373 VSS 0.28552f
C10479 a_46220_n6373 VSS 0.284099f
C10480 a_45772_n6373 VSS 0.284099f
C10481 a_45324_n6373 VSS 0.284099f
C10482 a_44876_n6373 VSS 0.285753f
C10483 a_44428_n6373 VSS 0.285466f
C10484 a_43980_n6373 VSS 0.285633f
C10485 a_43532_n6373 VSS 0.285633f
C10486 a_43084_n6373 VSS 0.288993f
C10487 a_42636_n6373 VSS 0.290707f
C10488 a_42188_n6373 VSS 0.292301f
C10489 a_41740_n6373 VSS 0.315404f
C10490 a_41292_n6373 VSS 0.299343f
C10491 a_40396_n6373 VSS 0.276502f
C10492 a_39948_n6373 VSS 0.293901f
C10493 a_39500_n6373 VSS 0.287277f
C10494 a_30740_n7464 VSS 0.538004f
C10495 a_31068_n6276 VSS 0.012971f
C10496 a_30616_n6221 VSS 0.281728f
C10497 a_30111_n6221 VSS 0.145471f
C10498 a_30808_n6334 VSS 0.335295f
C10499 a_30215_n6265 VSS 1.87623f
C10500 a_29123_n6679 VSS 1.7533f
C10501 a_30320_n6636 VSS 1.36638f
C10502 a_29559_n6456 VSS 0.37127f
C10503 a_29211_n6724 VSS 0.773786f
C10504 a_25972_n6276 VSS 1.78731f
C10505 a_25524_n6635 VSS 0.467668f
C10506 a_25612_n6679 VSS 1.74563f
C10507 a_24573_n6724 VSS 0.745589f
C10508 a_23949_n6724 VSS 0.730968f
C10509 a_21812_n6643 VSS 0.991711f
C10510 a_23619_n6724 VSS 0.612913f
C10511 a_22968_n6679 VSS 0.407973f
C10512 a_47900_n5940 VSS 0.300977f
C10513 a_47452_n5940 VSS 0.294024f
C10514 a_47004_n5940 VSS 0.29129f
C10515 a_46556_n5940 VSS 0.287668f
C10516 a_46108_n5940 VSS 0.285997f
C10517 a_45660_n5940 VSS 0.285997f
C10518 a_45212_n5940 VSS 0.289733f
C10519 a_47812_n5896 VSS 0.483823f
C10520 a_47364_n5896 VSS 0.46949f
C10521 a_46916_n5896 VSS 0.46798f
C10522 a_46468_n5896 VSS 0.461248f
C10523 a_46020_n5896 VSS 0.461248f
C10524 a_45572_n5896 VSS 0.461248f
C10525 a_45124_n5896 VSS 0.478762f
C10526 a_44204_n5940 VSS 0.271296f
C10527 a_43756_n5940 VSS 0.290733f
C10528 a_43308_n5940 VSS 0.291738f
C10529 a_42860_n5940 VSS 0.290233f
C10530 a_42412_n5940 VSS 0.292287f
C10531 a_41964_n5940 VSS 0.294993f
C10532 a_41516_n5940 VSS 0.325002f
C10533 a_41068_n5940 VSS 0.294181f
C10534 a_40620_n5940 VSS 0.291215f
C10535 a_40172_n5940 VSS 0.289616f
C10536 a_37820_n5940 VSS 0.243619f
C10537 a_37372_n5940 VSS 0.288635f
C10538 a_44116_n5896 VSS 0.483511f
C10539 a_43668_n5896 VSS 0.479297f
C10540 a_43220_n5896 VSS 0.472798f
C10541 a_42772_n5896 VSS 0.474227f
C10542 a_42324_n5896 VSS 0.476361f
C10543 a_41876_n5896 VSS 0.483976f
C10544 a_41428_n5896 VSS 0.492811f
C10545 a_40980_n5896 VSS 0.477147f
C10546 a_40532_n5896 VSS 0.460293f
C10547 a_40084_n5896 VSS 0.464922f
C10548 a_39357_n5364 VSS 0.775535f
C10549 a_38733_n5431 VSS 0.752879f
C10550 a_38403_n5503 VSS 0.621032f
C10551 a_37732_n5896 VSS 0.469875f
C10552 a_37284_n5896 VSS 0.480451f
C10553 a_29612_n8292 VSS 0.768578f
C10554 a_36773_n5468 VSS 0.59197f
C10555 a_22772_n5808 VSS 0.012971f
C10556 a_24128_n5408 VSS 0.145471f
C10557 a_23816_n5408 VSS 0.372165f
C10558 a_24233_n5548 VSS 0.768319f
C10559 a_22568_n5808 VSS 0.335295f
C10560 a_22364_n5808 VSS 0.075356f
C10561 a_22876_n5852 VSS 0.280902f
C10562 a_22264_n5852 VSS 0.417568f
C10563 a_22016_n5825 VSS 1.86844f
C10564 a_21604_n5412 VSS 1.46392f
C10565 a_47924_n4708 VSS 0.474295f
C10566 a_47476_n4708 VSS 0.461553f
C10567 a_47028_n4708 VSS 0.45987f
C10568 a_46580_n4708 VSS 0.457171f
C10569 a_46132_n4708 VSS 0.45666f
C10570 a_45684_n4708 VSS 0.45666f
C10571 a_45236_n4708 VSS 0.45666f
C10572 a_44788_n4708 VSS 0.471552f
C10573 a_44340_n4708 VSS 0.469522f
C10574 a_43892_n4708 VSS 0.470794f
C10575 a_43444_n4708 VSS 0.471552f
C10576 a_42996_n4708 VSS 0.474071f
C10577 a_42548_n4708 VSS 0.47587f
C10578 a_42100_n4708 VSS 0.47863f
C10579 a_41652_n4708 VSS 0.512838f
C10580 a_41204_n4708 VSS 0.493052f
C10581 a_40420_n4708 VSS 0.473086f
C10582 a_39972_n4708 VSS 0.4677f
C10583 a_39524_n4708 VSS 0.460411f
C10584 a_39076_n4708 VSS 0.474173f
C10585 a_38628_n4708 VSS 0.453101f
C10586 a_38180_n4708 VSS 0.476057f
C10587 a_48012_n4805 VSS 0.321039f
C10588 a_47564_n4805 VSS 0.290098f
C10589 a_47116_n4805 VSS 0.288045f
C10590 a_46668_n4805 VSS 0.28552f
C10591 a_46220_n4805 VSS 0.284099f
C10592 a_45772_n4805 VSS 0.284099f
C10593 a_45324_n4805 VSS 0.284099f
C10594 a_44876_n4805 VSS 0.285753f
C10595 a_44428_n4805 VSS 0.284269f
C10596 a_43980_n4805 VSS 0.284262f
C10597 a_43532_n4805 VSS 0.284262f
C10598 a_43084_n4805 VSS 0.287633f
C10599 a_42636_n4805 VSS 0.289347f
C10600 a_42188_n4805 VSS 0.2916f
C10601 a_41740_n4805 VSS 0.314382f
C10602 a_41292_n4805 VSS 0.298328f
C10603 a_40508_n4805 VSS 0.275489f
C10604 a_40060_n4805 VSS 0.288963f
C10605 a_39612_n4805 VSS 0.285404f
C10606 a_39164_n4805 VSS 0.284099f
C10607 a_38716_n4805 VSS 0.290116f
C10608 a_38268_n4805 VSS 0.289828f
C10609 a_28548_n5112 VSS 3.23851f
C10610 a_27414_n5112 VSS 0.683874f
C10611 a_27190_n5112 VSS 0.753243f
C10612 a_24180_n5112 VSS 0.507137f
C10613 a_22564_n5112 VSS 0.174573f
C10614 a_22220_n9860 VSS 0.796733f
C10615 a_23228_n6679 VSS 0.563535f
C10616 a_23207_n4708 VSS 0.026799f
C10617 a_26358_n4618 VSS 0.944967f
C10618 a_26154_n4536 VSS 0.744616f
C10619 a_25530_n5112 VSS 0.77599f
C10620 a_25237_n5895 VSS 0.840039f
C10621 a_24672_n11339 VSS 1.29625f
C10622 a_24492_n5156 VSS 1.57238f
C10623 a_23887_n5156 VSS 0.601378f
C10624 a_23479_n5156 VSS 1.43667f
C10625 a_22544_n4690 VSS 0.752934f
C10626 a_22444_n5156 VSS 3.90139f
C10627 a_21604_n5067 VSS 0.467968f
C10628 a_47900_n4372 VSS 0.300977f
C10629 a_47452_n4372 VSS 0.294024f
C10630 a_47004_n4372 VSS 0.29129f
C10631 a_46556_n4372 VSS 0.287668f
C10632 a_46108_n4372 VSS 0.285997f
C10633 a_45660_n4372 VSS 0.285997f
C10634 a_45212_n4372 VSS 0.289177f
C10635 a_47812_n4328 VSS 0.483823f
C10636 a_47364_n4328 VSS 0.46949f
C10637 a_46916_n4328 VSS 0.46798f
C10638 a_46468_n4328 VSS 0.461248f
C10639 a_46020_n4328 VSS 0.461248f
C10640 a_45572_n4328 VSS 0.461248f
C10641 a_45124_n4328 VSS 0.473068f
C10642 a_44540_n4372 VSS 0.291094f
C10643 a_44092_n4372 VSS 0.288363f
C10644 a_43644_n4372 VSS 0.286188f
C10645 a_43196_n4372 VSS 0.289237f
C10646 a_42748_n4372 VSS 0.290776f
C10647 a_42300_n4372 VSS 0.292239f
C10648 a_41852_n4372 VSS 0.299523f
C10649 a_41404_n4372 VSS 0.307822f
C10650 a_40956_n4372 VSS 0.293449f
C10651 a_40508_n4372 VSS 0.285951f
C10652 a_40060_n4372 VSS 0.284326f
C10653 a_39612_n4372 VSS 0.281201f
C10654 a_39164_n4372 VSS 0.281827f
C10655 a_33868_n4240 VSS 0.014304f
C10656 a_34736_n3840 VSS 0.081636f
C10657 a_44452_n4328 VSS 0.471915f
C10658 a_44004_n4328 VSS 0.461396f
C10659 a_43556_n4328 VSS 0.461394f
C10660 a_43108_n4328 VSS 0.464381f
C10661 a_42660_n4328 VSS 0.465992f
C10662 a_42212_n4328 VSS 0.4631f
C10663 a_41764_n4328 VSS 0.484654f
C10664 a_41316_n4328 VSS 0.465383f
C10665 a_40868_n4328 VSS 0.47782f
C10666 a_40420_n4328 VSS 0.459897f
C10667 a_39972_n4328 VSS 0.457363f
C10668 a_39524_n4328 VSS 0.455281f
C10669 a_39076_n4328 VSS 0.494165f
C10670 a_36520_n3868 VSS 0.457201f
C10671 a_35848_n3868 VSS 0.404802f
C10672 a_33416_n4240 VSS 0.283982f
C10673 a_28225_n4327 VSS 0.030139f
C10674 a_32911_n4240 VSS 0.145471f
C10675 a_33608_n4284 VSS 0.341237f
C10676 a_33015_n4284 VSS 1.87991f
C10677 a_33120_n3884 VSS 1.40024f
C10678 a_32359_n4372 VSS 0.32423f
C10679 a_31787_n3969 VSS 1.0515f
C10680 a_27540_n3797 VSS 0.438522f
C10681 a_28144_n4708 VSS 1.58022f
C10682 a_22772_n4240 VSS 0.012971f
C10683 a_24128_n3840 VSS 0.145471f
C10684 a_26271_n4306 VSS 0.619147f
C10685 a_26047_n4328 VSS 0.769961f
C10686 a_25423_n4328 VSS 0.724755f
C10687 a_23816_n3840 VSS 0.376201f
C10688 a_24233_n3980 VSS 0.764616f
C10689 a_22568_n4240 VSS 0.335295f
C10690 a_22364_n4240 VSS 0.075356f
C10691 a_22876_n4284 VSS 0.280882f
C10692 a_21792_n7464 VSS 0.655404f
C10693 a_22016_n4257 VSS 1.86962f
C10694 a_21604_n3844 VSS 1.42449f
C10695 a_47924_n3140 VSS 0.474295f
C10696 a_47476_n3140 VSS 0.461553f
C10697 a_47028_n3140 VSS 0.45987f
C10698 a_46580_n3140 VSS 0.457171f
C10699 a_46132_n3140 VSS 0.45666f
C10700 a_45684_n3140 VSS 0.45666f
C10701 a_45236_n3140 VSS 0.45666f
C10702 a_44788_n3140 VSS 0.471552f
C10703 a_44340_n3140 VSS 0.457943f
C10704 a_43892_n3140 VSS 0.457916f
C10705 a_43444_n3140 VSS 0.458675f
C10706 a_42996_n3140 VSS 0.461237f
C10707 a_42548_n3140 VSS 0.463036f
C10708 a_42100_n3140 VSS 0.465768f
C10709 a_41652_n3140 VSS 0.499298f
C10710 a_41204_n3140 VSS 0.482004f
C10711 a_40308_n3140 VSS 0.476847f
C10712 a_39860_n3140 VSS 0.467642f
C10713 a_39412_n3140 VSS 0.490122f
C10714 a_48012_n3237 VSS 0.32267f
C10715 a_47564_n3237 VSS 0.291728f
C10716 a_47116_n3237 VSS 0.289675f
C10717 a_46668_n3237 VSS 0.28715f
C10718 a_46220_n3237 VSS 0.285729f
C10719 a_45772_n3237 VSS 0.285729f
C10720 a_45324_n3237 VSS 0.285729f
C10721 a_44876_n3237 VSS 0.287383f
C10722 a_44428_n3237 VSS 0.285729f
C10723 a_43980_n3237 VSS 0.285729f
C10724 a_43532_n3237 VSS 0.285729f
C10725 a_43084_n3237 VSS 0.289162f
C10726 a_42636_n3237 VSS 0.290759f
C10727 a_42188_n3237 VSS 0.29171f
C10728 a_41740_n3237 VSS 0.314492f
C10729 a_41292_n3237 VSS 0.298352f
C10730 a_40396_n3237 VSS 0.274684f
C10731 a_39948_n3237 VSS 0.294015f
C10732 a_39500_n3237 VSS 0.287485f
C10733 a_37585_n3140 VSS 0.481235f
C10734 a_22052_n4708 VSS 3.03943f
C10735 a_36112_n3456 VSS 0.146447f
C10736 a_36217_n3500 VSS 0.772953f
C10737 a_35800_n3456 VSS 0.382017f
C10738 a_34756_n3140 VSS 0.025773f
C10739 a_34552_n3140 VSS 0.350062f
C10740 a_34348_n3140 VSS 0.077357f
C10741 a_34860_n3189 VSS 0.303448f
C10742 a_34000_n3140 VSS 1.88446f
C10743 a_29560_n3544 VSS 2.85239f
C10744 a_28583_n3140 VSS 0.027476f
C10745 a_33588_n3461 VSS 1.40594f
C10746 a_25600_n5895 VSS 1.21001f
C10747 a_27337_n3140 VSS 0.754186f
C10748 a_27932_n3543 VSS 0.72461f
C10749 a_27672_n3543 VSS 0.456931f
C10750 a_26607_n3544 VSS 0.635299f
C10751 a_26383_n2968 VSS 0.758526f
C10752 a_25759_n3544 VSS 0.76711f
C10753 a_25237_n4327 VSS 1.57171f
C10754 a_47900_n2804 VSS 0.300977f
C10755 a_47452_n2804 VSS 0.294024f
C10756 a_47004_n2804 VSS 0.29129f
C10757 a_46556_n2804 VSS 0.287668f
C10758 a_46108_n2804 VSS 0.285997f
C10759 a_45660_n2804 VSS 0.285997f
C10760 a_45212_n2804 VSS 0.289589f
C10761 a_47812_n2760 VSS 0.466214f
C10762 a_47364_n2760 VSS 0.451882f
C10763 a_46916_n2760 VSS 0.450371f
C10764 a_46468_n2760 VSS 0.443639f
C10765 a_46020_n2760 VSS 0.443639f
C10766 a_45572_n2760 VSS 0.443639f
C10767 a_45124_n2760 VSS 0.459814f
C10768 a_44316_n2804 VSS 0.271026f
C10769 a_43868_n2804 VSS 0.289079f
C10770 a_43420_n2804 VSS 0.285694f
C10771 a_42972_n2804 VSS 0.288461f
C10772 a_42524_n2804 VSS 0.290351f
C10773 a_42076_n2804 VSS 0.291794f
C10774 a_41628_n2804 VSS 0.328875f
C10775 a_41180_n2804 VSS 0.292742f
C10776 a_40732_n2804 VSS 0.293155f
C10777 a_37452_n3888 VSS 0.624379f
C10778 a_33188_n2672 VSS 0.014138f
C10779 a_44228_n2760 VSS 0.454391f
C10780 a_43780_n2760 VSS 0.438283f
C10781 a_43332_n2760 VSS 0.439994f
C10782 a_42884_n2760 VSS 0.453317f
C10783 a_42436_n2760 VSS 0.450996f
C10784 a_41988_n2760 VSS 0.459417f
C10785 a_41540_n2760 VSS 0.494166f
C10786 a_41092_n2760 VSS 0.462779f
C10787 a_40644_n2760 VSS 0.476662f
C10788 a_39357_n2228 VSS 0.735194f
C10789 a_38733_n2295 VSS 0.772075f
C10790 a_38403_n2367 VSS 0.63606f
C10791 a_34544_n2272 VSS 0.14937f
C10792 a_34232_n2272 VSS 0.336509f
C10793 a_34649_n2412 VSS 1.66785f
C10794 a_32984_n2672 VSS 0.337509f
C10795 a_32780_n2672 VSS 0.075356f
C10796 a_33292_n2716 VSS 0.29254f
C10797 a_32432_n2689 VSS 1.88297f
C10798 a_31392_n2760 VSS 0.435886f
C10799 a_31412_n2276 VSS 0.155702f
C10800 a_30555_n2729 VSS 0.541703f
C10801 a_27628_n3841 VSS 0.970421f
C10802 a_32020_n2276 VSS 1.38252f
C10803 a_31292_n2804 VSS 0.64044f
C10804 a_27348_n2672 VSS 0.071149f
C10805 a_28454_n2424 VSS 0.774455f
C10806 a_27452_n2716 VSS 0.497527f
C10807 a_25895_n2624 VSS 0.297033f
C10808 a_26499_n2732 VSS 0.344721f
C10809 a_23319_n2759 VSS 0.026799f
C10810 a_25139_n2704 VSS 0.049992f
C10811 a_25547_n2445 VSS 2.22501f
C10812 a_24771_n2804 VSS 1.59275f
C10813 a_23507_n2759 VSS 0.724379f
C10814 a_24403_n2414 VSS 0.672224f
C10815 a_22164_n2760 VSS 1.40173f
C10816 a_21716_n2229 VSS 0.462497f
C10817 a_22820_n2804 VSS 0.808028f
C10818 a_42116_n1976 VSS 0.010262f
C10819 a_47812_n1572 VSS 0.466214f
C10820 a_47364_n1572 VSS 0.451882f
C10821 a_46916_n1572 VSS 0.450371f
C10822 a_46468_n1572 VSS 0.438283f
C10823 a_46020_n1572 VSS 0.438283f
C10824 a_45572_n1572 VSS 0.438283f
C10825 a_45124_n1572 VSS 0.438283f
C10826 a_44676_n1572 VSS 0.469557f
C10827 a_44228_n1572 VSS 0.438283f
C10828 a_43780_n1572 VSS 0.438283f
C10829 a_43332_n1572 VSS 0.442252f
C10830 a_41204_n1572 VSS 0.48698f
C10831 a_34248_n3310 VSS 0.657613f
C10832 a_34953_n1572 VSS 0.568649f
C10833 a_32100_n1976 VSS 0.502431f
C10834 a_47900_n1669 VSS 0.299079f
C10835 a_47452_n1669 VSS 0.292126f
C10836 a_47004_n1669 VSS 0.289391f
C10837 a_46556_n1669 VSS 0.285046f
C10838 a_46108_n1669 VSS 0.281201f
C10839 a_45660_n1669 VSS 0.281201f
C10840 a_45212_n1669 VSS 0.281201f
C10841 a_44764_n1669 VSS 0.285973f
C10842 a_44316_n1669 VSS 0.281201f
C10843 a_43868_n1669 VSS 0.282953f
C10844 a_43420_n1669 VSS 0.287725f
C10845 a_42244_n1572 VSS 1.03701f
C10846 a_41684_n1976 VSS 0.461208f
C10847 a_41292_n1669 VSS 0.250124f
C10848 a_40196_n1884 VSS 0.363611f
C10849 a_37221_n3543 VSS 1.4205f
C10850 a_39648_n2020 VSS 0.354308f
C10851 a_38984_n1975 VSS 0.412169f
C10852 a_38312_n1975 VSS 0.414622f
C10853 a_37632_n2020 VSS 0.357515f
C10854 a_36388_n1572 VSS 1.1714f
C10855 a_36744_n1954 VSS 0.679566f
C10856 a_35940_n1931 VSS 0.424465f
C10857 a_35288_n1975 VSS 0.426362f
C10858 a_34223_n1976 VSS 0.643695f
C10859 a_33999_n1400 VSS 0.743696f
C10860 a_32308_n1976 VSS 0.595282f
C10861 a_33375_n1976 VSS 0.752979f
C10862 a_32860_n2020 VSS 0.687231f
C10863 a_32636_n2020 VSS 0.613231f
C10864 a_31348_n1931 VSS 0.407668f
C10865 a_27988_n4328 VSS 5.12978f
C10866 a_30584_n1954 VSS 0.665481f
C10867 a_29519_n1976 VSS 0.631196f
C10868 a_29295_n1400 VSS 0.753601f
C10869 a_28671_n1976 VSS 0.746594f
C10870 a_26495_n1976 VSS 0.630748f
C10871 a_26271_n1400 VSS 0.760255f
C10872 a_25647_n1976 VSS 0.750217f
C10873 a_24315_n2759 VSS 0.807984f
C10874 a_24578_n2020 VSS 0.772101f
C10875 a_23954_n2020 VSS 0.741312f
C10876 a_23542_n1754 VSS 0.930509f
C10877 a_22918_n2020 VSS 0.737007f
C10878 a_22588_n2020 VSS 0.641847f
C10879 a_21828_n1931 VSS 0.455406f
C10880 a_21916_n1975 VSS 1.11175f
C10881 a_47900_n1236 VSS 0.299079f
C10882 a_47452_n1236 VSS 0.292126f
C10883 a_47004_n1236 VSS 0.289391f
C10884 a_46556_n1236 VSS 0.285769f
C10885 a_46108_n1236 VSS 0.284099f
C10886 a_45660_n1236 VSS 0.284099f
C10887 a_45212_n1236 VSS 0.287691f
C10888 a_47812_n1192 VSS 0.485254f
C10889 a_47364_n1192 VSS 0.470495f
C10890 a_46916_n1192 VSS 0.469363f
C10891 a_46468_n1192 VSS 0.461487f
C10892 a_46020_n1192 VSS 0.462614f
C10893 a_45572_n1192 VSS 0.461264f
C10894 a_45124_n1192 VSS 0.477439f
C10895 a_44316_n1236 VSS 0.267773f
C10896 a_43556_n661 VSS 0.419665f
C10897 a_42972_n1236 VSS 0.250152f
C10898 a_44228_n1192 VSS 0.491623f
C10899 a_42884_n1192 VSS 0.479828f
C10900 a_42157_n660 VSS 0.789429f
C10901 a_41533_n727 VSS 0.817043f
C10902 a_41203_n799 VSS 0.691696f
C10903 a_39357_n660 VSS 0.721727f
C10904 a_38733_n727 VSS 0.763322f
C10905 a_38403_n799 VSS 0.63667f
C10906 a_33077_n1191 VSS 0.638418f
C10907 a_30612_n1104 VSS 0.012971f
C10908 a_31968_n704 VSS 0.145471f
C10909 a_35119_n1170 VSS 0.627756f
C10910 a_34895_n1192 VSS 0.789274f
C10911 a_34271_n1192 VSS 0.761513f
C10912 a_33252_n1192 VSS 0.68216f
C10913 a_31656_n704 VSS 0.38384f
C10914 a_32073_n844 VSS 0.766357f
C10915 a_30408_n1104 VSS 0.335295f
C10916 a_30204_n1104 VSS 0.075356f
C10917 a_30716_n1148 VSS 0.283145f
C10918 a_29856_n1121 VSS 1.87444f
C10919 a_29444_n708 VSS 1.47747f
C10920 a_25524_n708 VSS 0.150169f
C10921 a_22772_n1104 VSS 0.012971f
C10922 a_24128_n704 VSS 0.145471f
C10923 a_27279_n1170 VSS 0.643831f
C10924 a_27055_n1192 VSS 0.739245f
C10925 a_26431_n1192 VSS 0.724282f
C10926 a_23816_n704 VSS 0.37752f
C10927 a_24233_n844 VSS 0.771709f
C10928 a_22568_n1104 VSS 0.335295f
C10929 a_22364_n1104 VSS 0.075356f
C10930 a_22876_n1148 VSS 0.280882f
C10931 a_22016_n1121 VSS 1.86843f
C10932 a_21604_n708 VSS 1.43206f
C10933 a_47924_n4 VSS 0.48572f
C10934 a_47476_n4 VSS 0.470088f
C10935 a_47028_n4 VSS 0.468405f
C10936 a_46580_n4 VSS 0.461869f
C10937 a_46132_n4 VSS 0.461358f
C10938 a_45684_n4 VSS 0.461358f
C10939 a_45236_n4 VSS 0.467456f
C10940 a_48012_n101 VSS 0.320457f
C10941 a_47564_n101 VSS 0.29448f
C10942 a_47116_n101 VSS 0.291209f
C10943 a_46668_n101 VSS 0.286979f
C10944 a_46220_n101 VSS 0.286275f
C10945 a_45772_n101 VSS 0.286328f
C10946 a_45324_n101 VSS 0.287579f
C10947 a_42948_n1976 VSS 0.940171f
C10948 a_44509_n452 VSS 0.778838f
C10949 a_43885_n452 VSS 0.761713f
C10950 a_42772_n4 VSS 0.470239f
C10951 a_42324_n4 VSS 0.489014f
C10952 a_43555_n452 VSS 0.630853f
C10953 a_42860_n101 VSS 0.255314f
C10954 a_42412_n101 VSS 0.295529f
C10955 a_41336_n407 VSS 0.463155f
C10956 a_39556_n4 VSS 1.05102f
C10957 a_38996_n408 VSS 0.408723f
C10958 a_39308_n452 VSS 0.773468f
C10959 a_33940_n408 VSS 0.010308f
C10960 a_37680_n320 VSS 0.145471f
C10961 a_37785_n364 VSS 0.760252f
C10962 a_37368_n320 VSS 0.381668f
C10963 a_36324_n4 VSS 0.013806f
C10964 a_36120_n4 VSS 0.336978f
C10965 a_35916_n4 VSS 0.076765f
C10966 a_36428_n53 VSS 0.291418f
C10967 a_35568_n4 VSS 1.88155f
C10968 a_35156_n325 VSS 1.44197f
C10969 a_34068_n4 VSS 1.05472f
C10970 a_33508_n408 VSS 0.474895f
C10971 a_32262_n452 VSS 0.739063f
C10972 a_31405_n452 VSS 0.716235f
C10973 a_30781_n452 VSS 0.746299f
C10974 a_28352_n320 VSS 0.078257f
C10975 a_30451_n452 VSS 0.630544f
C10976 a_28456_n364 VSS 0.43337f
C10977 a_27484_n4 VSS 0.021364f
C10978 a_27032_51 VSS 0.292581f
C10979 a_26527_51 VSS 0.146012f
C10980 a_27224_n62 VSS 0.365646f
C10981 a_26631_7 VSS 1.90045f
C10982 a_26736_n364 VSS 1.47868f
C10983 a_25975_n184 VSS 0.379121f
C10984 a_25627_n452 VSS 0.756937f
C10985 a_24628_n363 VSS 0.439973f
C10986 a_48012_332 VSS 0.320484f
C10987 a_42604_n2020 VSS 0.813398f
C10988 a_45660_332 VSS 0.245521f
C10989 a_45212_332 VSS 0.290598f
C10990 a_47924_376 VSS 0.487939f
C10991 a_47197_908 VSS 0.773094f
C10992 a_46573_841 VSS 0.761702f
C10993 a_46243_769 VSS 0.617704f
C10994 a_45572_376 VSS 0.463102f
C10995 a_45124_376 VSS 0.476517f
C10996 a_44540_332 VSS 0.287751f
C10997 a_39804_464 VSS 0.013617f
C10998 a_40672_864 VSS 0.076736f
C10999 a_44452_376 VSS 0.487674f
C11000 a_40260_n408 VSS 0.932446f
C11001 a_43725_908 VSS 0.745642f
C11002 a_43101_841 VSS 0.742423f
C11003 a_42771_769 VSS 0.624525f
C11004 a_40776_770 VSS 0.554823f
C11005 a_39352_464 VSS 0.281325f
C11006 a_38847_464 VSS 0.145471f
C11007 a_39544_420 VSS 0.336662f
C11008 a_38951_420 VSS 1.8731f
C11009 a_39056_820 VSS 1.46131f
C11010 a_38295_332 VSS 0.376634f
C11011 a_37947_332 VSS 0.766436f
C11012 a_30104_n1148 VSS 0.846189f
C11013 a_35816_n174 VSS 0.422378f
C11014 a_31076_376 VSS 0.771632f
C11015 a_35119_398 VSS 0.638006f
C11016 a_34895_376 VSS 0.769933f
C11017 a_34271_376 VSS 0.722131f
C11018 a_34403_332 VSS 0.70477f
C11019 a_33533_908 VSS 0.738472f
C11020 a_32909_841 VSS 0.769174f
C11021 a_32579_769 VSS 0.632739f
C11022 a_24631_n3588 VSS 2.09046f
C11023 a_30372_376 VSS 1.00216f
C11024 a_29812_860 VSS 0.457491f
C11025 a_28004_860 VSS 0.013868f
C11026 a_23004_n2332 VSS 0.807356f
C11027 a_28132_376 VSS 1.06548f
C11028 a_28492_332 VSS 0.744388f
C11029 a_27572_860 VSS 0.441377f
C11030 a_25817_804 VSS 0.658691f
C11031 a_25137_864 VSS 0.049992f
C11032 a_24913_864 VSS 1.58883f
C11033 a_23524_464 VSS 0.069774f
C11034 a_23728_464 VSS 0.341193f
C11035 a_24041_816 VSS 0.296309f
C11036 a_23404_816 VSS 0.57714f
C11037 a_23136_447 VSS 2.24028f
C11038 a_22116_860 VSS 0.155702f
C11039 a_45012_1564 VSS 0.468181f
C11040 a_43644_n705 VSS 1.90165f
C11041 a_40652_n1572 VSS 2.57262f
C11042 a_45100_1467 VSS 0.267097f
C11043 a_43728_1248 VSS 0.145471f
C11044 a_43833_1204 VSS 0.766457f
C11045 a_43416_1248 VSS 0.390893f
C11046 a_42372_1564 VSS 0.01607f
C11047 a_42168_1564 VSS 0.34284f
C11048 a_41964_1564 VSS 0.080241f
C11049 a_42476_1515 VSS 0.294665f
C11050 a_41864_1394 VSS 0.911277f
C11051 a_41616_1564 VSS 1.91592f
C11052 a_36192_1248 VSS 0.076553f
C11053 a_41204_1243 VSS 1.48923f
C11054 a_37844_1564 VSS 1.42386f
C11055 a_37396_1205 VSS 0.43769f
C11056 a_35849_n1192 VSS 0.738216f
C11057 a_35324_1564 VSS 0.017071f
C11058 a_34872_1619 VSS 0.313786f
C11059 a_34367_1619 VSS 0.149048f
C11060 a_35064_1506 VSS 0.347616f
C11061 a_34471_1575 VSS 1.91194f
C11062 a_34576_1204 VSS 1.47335f
C11063 a_33815_1384 VSS 0.398776f
C11064 a_33467_1116 VSS 0.770252f
C11065 a_31856_1248 VSS 0.145471f
C11066 a_31961_1204 VSS 0.770545f
C11067 a_31544_1248 VSS 0.380574f
C11068 a_30500_1564 VSS 0.012971f
C11069 a_30296_1564 VSS 0.335295f
C11070 a_30092_1564 VSS 0.075356f
C11071 a_30604_1515 VSS 0.28372f
C11072 a_28836_376 VSS 0.66489f
C11073 a_29744_1564 VSS 1.87261f
C11074 a_29332_1243 VSS 1.38012f
C11075 a_28048_1248 VSS 0.167341f
C11076 a_28153_1204 VSS 0.78733f
C11077 a_27736_1248 VSS 0.389684f
C11078 a_26692_1564 VSS 0.013972f
C11079 a_26488_1564 VSS 0.339707f
C11080 a_26284_1564 VSS 0.075395f
C11081 a_26796_1515 VSS 0.289509f
C11082 a_22096_376 VSS 0.653679f
C11083 a_25936_1564 VSS 1.89505f
C11084 a_25524_1243 VSS 1.46152f
C11085 a_24628_1252 VSS 0.352188f
C11086 a_47452_1900 VSS 0.2873f
C11087 a_47364_1944 VSS 0.510532f
C11088 a_44004_n1192 VSS 1.88665f
C11089 a_40196_1944 VSS 2.76982f
C11090 a_39748_2475 VSS 0.444153f
C11091 a_37859_377 VSS 1.86759f
C11092 a_36388_1944 VSS 1.63678f
C11093 a_35940_2475 VSS 0.448246f
C11094 a_25084_1564 VSS 1.65327f
C11095 a_31324_n4372 VSS 1.42389f
C11096 a_28736_1944 VSS 0.690581f
C11097 a_22500_n1976 VSS 1.46785f
C11098 a_32132_2428 VSS 0.369821f
C11099 a_26607_1966 VSS 0.646483f
C11100 a_26383_1944 VSS 0.784286f
C11101 a_25759_1944 VSS 0.775391f
C11102 a_22052_1944 VSS 2.61803f
C11103 a_21604_2475 VSS 0.484046f
C11104 a_21692_2431 VSS 1.50437f
C11105 a_n199_2852 VSS 3.53357f
C11106 a_7119_4292 VSS 1.95081f
C11107 a_3025_2852 VSS 1.99373f
C11108 a_137_4292 VSS 2.97928f
C11109 a_21692_n7508.t0 VSS 0.051698f
C11110 a_21692_n7508.t3 VSS 0.084306f
C11111 a_21692_n7508.t2 VSS 0.155014f
C11112 a_21692_n7508.n0 VSS 2.02125f
C11113 a_21692_n7508.n1 VSS 3.04327f
C11114 a_21692_n7508.t1 VSS 0.144462f
C11115 a_27225_n1572.t1 VSS 3.21439f
C11116 a_27225_n1572.t2 VSS 0.129716f
C11117 a_27225_n1572.t3 VSS 0.100898f
C11118 a_27225_n1572.n0 VSS 2.67166f
C11119 a_27225_n1572.t0 VSS 0.083341f
C11120 a_24716_1208.t1 VSS 0.203488f
C11121 a_24716_1208.t0 VSS 0.032437f
C11122 a_24716_1208.t4 VSS 0.025467f
C11123 a_24716_1208.t5 VSS 0.051544f
C11124 a_24716_1208.n0 VSS 0.168073f
C11125 a_24716_1208.t2 VSS 0.040977f
C11126 a_24716_1208.t3 VSS 0.026094f
C11127 a_24716_1208.n1 VSS 0.434344f
C11128 a_24716_1208.n2 VSS 1.21757f
C11129 a_22668_n14864.t0 VSS 0.024858f
C11130 a_22668_n14864.t3 VSS 0.040536f
C11131 a_22668_n14864.t2 VSS 0.074535f
C11132 a_22668_n14864.n0 VSS 0.817562f
C11133 a_22668_n14864.n1 VSS 1.37305f
C11134 a_22668_n14864.t1 VSS 0.069461f
C11135 a_25795_n2716.t1 VSS 0.421531f
C11136 a_25795_n2716.t0 VSS 0.038068f
C11137 a_25795_n2716.t4 VSS 0.175684f
C11138 a_25795_n2716.t5 VSS 0.231525f
C11139 a_25795_n2716.t3 VSS 0.13409f
C11140 a_25795_n2716.t2 VSS 0.450407f
C11141 a_25795_n2716.t7 VSS 0.539579f
C11142 a_25795_n2716.t6 VSS 0.293265f
C11143 a_25795_n2716.n0 VSS 0.115851f
C11144 a_22276_n1572.t1 VSS 11.2686f
C11145 a_22276_n1572.t0 VSS 0.087018f
C11146 a_22276_n1572.t2 VSS 0.25315f
C11147 a_22276_n1572.t3 VSS 0.133353f
C11148 a_22276_n1572.n0 VSS 9.05784f
C11149 a_33820_n452.t1 VSS 1.55001f
C11150 a_33820_n452.t3 VSS 0.127918f
C11151 a_33820_n452.t2 VSS 0.074361f
C11152 a_33820_n452.n0 VSS 0.875361f
C11153 a_33820_n452.t0 VSS 0.072355f
C11154 a_24731_n3124.t0 VSS 1.01565f
C11155 a_24731_n3124.t1 VSS 0.022888f
C11156 a_24731_n3124.t5 VSS 0.029649f
C11157 a_24731_n3124.t3 VSS 0.034279f
C11158 a_24731_n3124.n0 VSS 0.102687f
C11159 a_24731_n3124.t4 VSS 0.029649f
C11160 a_24731_n3124.t2 VSS 0.034279f
C11161 a_24731_n3124.n1 VSS 0.192025f
C11162 a_24731_n3124.n2 VSS 1.73889f
C11163 a_27001_n4328.t1 VSS 1.19113f
C11164 a_27001_n4328.t2 VSS 0.025396f
C11165 a_27001_n4328.t3 VSS 0.046696f
C11166 a_27001_n4328.n0 VSS 0.80663f
C11167 a_27001_n4328.t0 VSS 0.030153f
C11168 a_25539_n407.t1 VSS 0.124689f
C11169 a_25539_n407.t2 VSS 0.031355f
C11170 a_25539_n407.t4 VSS 0.016517f
C11171 a_25539_n407.n0 VSS 0.535105f
C11172 a_25539_n407.t3 VSS 0.015176f
C11173 a_25539_n407.t5 VSS 0.030715f
C11174 a_25539_n407.n1 VSS 0.145872f
C11175 a_25539_n407.n2 VSS 1.17941f
C11176 a_25539_n407.t0 VSS 0.021158f
C11177 a_23999_n2320.t1 VSS 0.196386f
C11178 a_23999_n2320.n0 VSS 1.45648f
C11179 a_23999_n2320.t0 VSS 0.027124f
C11180 a_23999_n2320.t6 VSS 0.040197f
C11181 a_23999_n2320.t2 VSS 0.021175f
C11182 a_23999_n2320.n1 VSS 0.533932f
C11183 a_23999_n2320.t5 VSS 0.039376f
C11184 a_23999_n2320.t7 VSS 0.019455f
C11185 a_23999_n2320.n2 VSS 0.106985f
C11186 a_23999_n2320.t4 VSS 0.038875f
C11187 a_23999_n2320.t3 VSS 0.0363f
C11188 a_23999_n2320.n3 VSS 0.083714f
C11189 a_29263_n3588.n0 VSS 2.27936f
C11190 a_29263_n3588.t0 VSS 0.135931f
C11191 a_29263_n3588.t1 VSS 0.076605f
C11192 a_29263_n3588.t3 VSS 0.113362f
C11193 a_29263_n3588.t2 VSS 0.120716f
C11194 a_29263_n3588.n1 VSS 1.47402f
C11195 a_23703_n5156.t0 VSS 0.026938f
C11196 a_23703_n5156.t1 VSS 0.046225f
C11197 a_23703_n5156.t5 VSS 0.023961f
C11198 a_23703_n5156.t6 VSS 0.029703f
C11199 a_23703_n5156.n0 VSS 0.053571f
C11200 a_23703_n5156.t4 VSS 0.023961f
C11201 a_23703_n5156.t7 VSS 0.029703f
C11202 a_23703_n5156.n1 VSS 0.044893f
C11203 a_23703_n5156.t2 VSS 0.029776f
C11204 a_23703_n5156.t3 VSS 0.023878f
C11205 a_23703_n5156.n2 VSS 0.044056f
C11206 a_23703_n5156.t9 VSS 0.029776f
C11207 a_23703_n5156.t11 VSS 0.023878f
C11208 a_23703_n5156.n3 VSS 0.055439f
C11209 a_23703_n5156.n4 VSS 0.403288f
C11210 a_23703_n5156.t8 VSS 0.029776f
C11211 a_23703_n5156.t10 VSS 0.023878f
C11212 a_23703_n5156.n5 VSS 0.044056f
C11213 a_23703_n5156.n6 VSS 0.583419f
C11214 a_23703_n5156.n7 VSS 0.333313f
C11215 a_23703_n5156.n8 VSS 0.318558f
C11216 a_23703_n5156.n9 VSS 0.07795f
C11217 a_26172_n14564.t0 VSS 1.88846f
C11218 a_26172_n14564.t1 VSS 0.046908f
C11219 a_26172_n14564.t2 VSS 0.060647f
C11220 a_26172_n14564.t3 VSS 0.050506f
C11221 a_26172_n14564.n0 VSS 1.25348f
C11222 a_28940_n2406.n0 VSS 0.484896f
C11223 a_28940_n2406.t1 VSS 0.072946f
C11224 a_28940_n2406.t0 VSS 0.046918f
C11225 a_28940_n2406.t4 VSS 0.061123f
C11226 a_28940_n2406.t5 VSS 0.075768f
C11227 a_28940_n2406.n1 VSS 0.136126f
C11228 a_28940_n2406.t6 VSS 0.061123f
C11229 a_28940_n2406.t7 VSS 0.075768f
C11230 a_28940_n2406.n2 VSS 0.217979f
C11231 a_28940_n2406.n3 VSS 1.34071f
C11232 a_28940_n2406.t3 VSS 0.064299f
C11233 a_28940_n2406.t2 VSS 0.07342f
C11234 a_28940_n2406.n4 VSS 0.299869f
C11235 a_28940_n2406.n5 VSS 2.18905f
C11236 a_22892_n5156.t0 VSS 0.077901f
C11237 a_22892_n5156.t2 VSS 0.014468f
C11238 a_22892_n5156.t1 VSS 0.047364f
C11239 a_22892_n5156.t4 VSS 0.059049f
C11240 a_22892_n5156.t3 VSS 0.04805f
C11241 a_22892_n5156.n0 VSS 0.809735f
C11242 a_22892_n5156.n1 VSS 1.14343f
C11243 a_25076_n4.t0 VSS 0.048052f
C11244 a_25076_n4.t3 VSS 0.129528f
C11245 a_25076_n4.t2 VSS 0.1269f
C11246 a_25076_n4.n0 VSS 3.06499f
C11247 a_25076_n4.n1 VSS 4.19625f
C11248 a_25076_n4.t1 VSS 0.134274f
C11249 a_28852_n8292.n0 VSS 1.11641f
C11250 a_28852_n8292.t0 VSS 0.076872f
C11251 a_28852_n8292.t1 VSS 0.043322f
C11252 a_28852_n8292.t3 VSS 0.067406f
C11253 a_28852_n8292.t2 VSS 0.061111f
C11254 a_28852_n8292.n1 VSS 0.734881f
C11255 a_29900_n10600.t1 VSS 0.353308f
C11256 a_29900_n10600.n0 VSS 0.100377f
C11257 a_29900_n10600.n1 VSS 0.056798f
C11258 a_29900_n10600.n2 VSS 0.09913f
C11259 a_29900_n10600.n3 VSS 2.37239f
C11260 a_29900_n10600.t0 VSS 0.042197f
C11261 a_29900_n10600.t8 VSS 0.055706f
C11262 a_29900_n10600.t5 VSS 0.064027f
C11263 a_29900_n10600.n4 VSS 0.397747f
C11264 a_29900_n10600.t2 VSS 0.054455f
C11265 a_29900_n10600.t3 VSS 0.070008f
C11266 a_29900_n10600.n5 VSS 0.50548f
C11267 a_29900_n10600.t7 VSS 0.04629f
C11268 a_29900_n10600.t6 VSS 0.04629f
C11269 a_29900_n10600.t9 VSS 0.067897f
C11270 a_29900_n10600.t4 VSS 0.067897f
C11271 a_23564_n3588.t1 VSS 3.32252f
C11272 a_23564_n3588.n0 VSS 0.181077f
C11273 a_23564_n3588.t0 VSS 0.03462f
C11274 a_23564_n3588.t8 VSS 0.097577f
C11275 a_23564_n3588.t7 VSS 0.090028f
C11276 a_23564_n3588.n1 VSS 0.149197f
C11277 a_23564_n3588.t9 VSS 0.097577f
C11278 a_23564_n3588.t3 VSS 0.101201f
C11279 a_23564_n3588.t2 VSS 0.085403f
C11280 a_23564_n3588.n2 VSS 0.158214f
C11281 a_23564_n3588.t4 VSS 0.085403f
C11282 a_23564_n3588.t6 VSS 0.097577f
C11283 a_23564_n3588.t5 VSS 0.090028f
C11284 a_23564_n3588.n3 VSS 3.10958f
C11285 a_34428_n452.t1 VSS 0.308462f
C11286 a_34428_n452.t5 VSS 0.084727f
C11287 a_34428_n452.t2 VSS 0.07103f
C11288 a_34428_n452.n0 VSS 0.348272f
C11289 a_34428_n452.t4 VSS 0.084069f
C11290 a_34428_n452.t7 VSS 0.044286f
C11291 a_34428_n452.n1 VSS 0.229272f
C11292 a_34428_n452.n2 VSS 1.24053f
C11293 a_34428_n452.t6 VSS 0.04069f
C11294 a_34428_n452.t3 VSS 0.082353f
C11295 a_34428_n452.n3 VSS 0.58424f
C11296 a_34428_n452.n4 VSS 1.02534f
C11297 a_34428_n452.t0 VSS 0.056728f
C11298 a_22264_n1148.t1 VSS 2.25706f
C11299 a_22264_n1148.t0 VSS 0.02328f
C11300 a_22264_n1148.t3 VSS 0.041214f
C11301 a_22264_n1148.t2 VSS 0.037836f
C11302 a_22264_n1148.n0 VSS 1.94061f
C11303 OUT[4].t3 VSS 0.016743f
C11304 OUT[4].t7 VSS 0.016743f
C11305 OUT[4].n0 VSS 0.033602f
C11306 OUT[4].t6 VSS 0.016743f
C11307 OUT[4].t0 VSS 0.016743f
C11308 OUT[4].n1 VSS 0.033602f
C11309 OUT[4].t5 VSS 0.016743f
C11310 OUT[4].t2 VSS 0.016743f
C11311 OUT[4].n2 VSS 0.040268f
C11312 OUT[4].n3 VSS 0.183905f
C11313 OUT[4].t11 VSS 0.034491f
C11314 OUT[4].t15 VSS 0.024911f
C11315 OUT[4].n4 VSS 0.060147f
C11316 OUT[4].t12 VSS 0.024911f
C11317 OUT[4].t9 VSS 0.034491f
C11318 OUT[4].n5 VSS 0.075016f
C11319 OUT[4].n6 VSS 0.188721f
C11320 OUT[4].t14 VSS 0.034491f
C11321 OUT[4].t8 VSS 0.024911f
C11322 OUT[4].n7 VSS 0.060147f
C11323 OUT[4].t13 VSS 0.034491f
C11324 OUT[4].t10 VSS 0.024911f
C11325 OUT[4].n8 VSS 0.076086f
C11326 OUT[4].n9 VSS 0.192426f
C11327 OUT[4].n10 VSS 0.147892f
C11328 OUT[4].n11 VSS 0.147892f
C11329 OUT[4].n12 VSS 0.105491f
C11330 OUT[4].t4 VSS 0.016743f
C11331 OUT[4].t1 VSS 0.016743f
C11332 OUT[4].n13 VSS 0.033486f
C11333 OUT[4].n14 VSS 0.303027f
C11334 a_27337_1944.t1 VSS 1.42714f
C11335 a_27337_1944.t2 VSS 0.053963f
C11336 a_27337_1944.t3 VSS 0.029348f
C11337 a_27337_1944.n0 VSS 1.1547f
C11338 a_27337_1944.t0 VSS 0.034846f
C11339 a_25836_n1236.n0 VSS 0.861143f
C11340 a_25836_n1236.n1 VSS 0.413711f
C11341 a_25836_n1236.n2 VSS 0.368431f
C11342 a_25836_n1236.n3 VSS 1.18288f
C11343 a_25836_n1236.t5 VSS 0.029835f
C11344 a_25836_n1236.t6 VSS 0.029835f
C11345 a_25836_n1236.t4 VSS 0.029835f
C11346 a_25836_n1236.n4 VSS 0.086493f
C11347 a_25836_n1236.t1 VSS 0.020013f
C11348 a_25836_n1236.t3 VSS 0.020013f
C11349 a_25836_n1236.n5 VSS 0.04514f
C11350 a_25836_n1236.t0 VSS 0.020013f
C11351 a_25836_n1236.t2 VSS 0.020013f
C11352 a_25836_n1236.n6 VSS 0.040161f
C11353 a_25836_n1236.t11 VSS 0.062159f
C11354 a_25836_n1236.t23 VSS 0.100113f
C11355 a_25836_n1236.n7 VSS 0.14612f
C11356 a_25836_n1236.t15 VSS 0.062159f
C11357 a_25836_n1236.t32 VSS 0.100113f
C11358 a_25836_n1236.n8 VSS 0.118799f
C11359 a_25836_n1236.n9 VSS 0.339414f
C11360 a_25836_n1236.t40 VSS 0.050852f
C11361 a_25836_n1236.t22 VSS 0.093501f
C11362 a_25836_n1236.n10 VSS 0.522937f
C11363 a_25836_n1236.t30 VSS 0.075793f
C11364 a_25836_n1236.t28 VSS 0.091049f
C11365 a_25836_n1236.n11 VSS 0.122119f
C11366 a_25836_n1236.t38 VSS 0.075793f
C11367 a_25836_n1236.t26 VSS 0.091049f
C11368 a_25836_n1236.n12 VSS 0.124494f
C11369 a_25836_n1236.t35 VSS 0.075793f
C11370 a_25836_n1236.t18 VSS 0.085574f
C11371 a_25836_n1236.t12 VSS 0.075793f
C11372 a_25836_n1236.n13 VSS 0.06139f
C11373 a_25836_n1236.t24 VSS 0.085574f
C11374 a_25836_n1236.n14 VSS 0.06961f
C11375 a_25836_n1236.n15 VSS 0.06961f
C11376 a_25836_n1236.n16 VSS 0.06139f
C11377 a_25836_n1236.t14 VSS 0.076784f
C11378 a_25836_n1236.t10 VSS 0.094362f
C11379 a_25836_n1236.n17 VSS 0.234277f
C11380 a_25836_n1236.t29 VSS 0.087933f
C11381 a_25836_n1236.t9 VSS 0.074376f
C11382 a_25836_n1236.n18 VSS 0.287904f
C11383 a_25836_n1236.n19 VSS 0.966277f
C11384 a_25836_n1236.t17 VSS 0.097279f
C11385 a_25836_n1236.t34 VSS 0.057714f
C11386 a_25836_n1236.n20 VSS 0.104825f
C11387 a_25836_n1236.n21 VSS 0.571311f
C11388 a_25836_n1236.t19 VSS 0.064784f
C11389 a_25836_n1236.t13 VSS 0.086418f
C11390 a_25836_n1236.n22 VSS 0.166468f
C11391 a_25836_n1236.n23 VSS 0.988864f
C11392 a_25836_n1236.n24 VSS 0.410401f
C11393 a_25836_n1236.t33 VSS 0.060917f
C11394 a_25836_n1236.n25 VSS 0.064303f
C11395 a_25836_n1236.t8 VSS 0.083309f
C11396 a_25836_n1236.n26 VSS 0.095533f
C11397 a_25836_n1236.t36 VSS 0.084057f
C11398 a_25836_n1236.n27 VSS 0.088741f
C11399 a_25836_n1236.t21 VSS 0.062472f
C11400 a_25836_n1236.n28 VSS 0.057096f
C11401 a_25836_n1236.t27 VSS 0.062472f
C11402 a_25836_n1236.n29 VSS 0.058791f
C11403 a_25836_n1236.t39 VSS 0.083309f
C11404 a_25836_n1236.t37 VSS 0.084057f
C11405 a_25836_n1236.n30 VSS 0.088741f
C11406 a_25836_n1236.n31 VSS 0.095533f
C11407 a_25836_n1236.t31 VSS 0.060917f
C11408 a_25836_n1236.n32 VSS 0.062618f
C11409 a_25836_n1236.n33 VSS 0.748332f
C11410 a_25836_n1236.t16 VSS 0.073432f
C11411 a_25836_n1236.t25 VSS 0.094593f
C11412 a_25836_n1236.n34 VSS 0.1324f
C11413 a_25836_n1236.t41 VSS 0.079613f
C11414 a_25836_n1236.t20 VSS 0.092533f
C11415 a_25836_n1236.n35 VSS 0.081762f
C11416 a_25836_n1236.n36 VSS 0.266934f
C11417 a_25836_n1236.n37 VSS 0.94934f
C11418 a_25836_n1236.n38 VSS 0.059671f
C11419 a_25836_n1236.t7 VSS 0.029835f
C11420 a_25019_n3588.t1 VSS 0.470585f
C11421 a_25019_n3588.n0 VSS 0.086187f
C11422 a_25019_n3588.n1 VSS 0.222166f
C11423 a_25019_n3588.n2 VSS 0.085598f
C11424 a_25019_n3588.t0 VSS 0.036503f
C11425 a_25019_n3588.t6 VSS 0.055539f
C11426 a_25019_n3588.t4 VSS 0.048189f
C11427 a_25019_n3588.n3 VSS 0.40702f
C11428 a_25019_n3588.t8 VSS 0.049483f
C11429 a_25019_n3588.t7 VSS 0.060811f
C11430 a_25019_n3588.n4 VSS 0.12062f
C11431 a_25019_n3588.n5 VSS 1.38305f
C11432 a_25019_n3588.t3 VSS 0.040077f
C11433 a_25019_n3588.t5 VSS 0.058887f
C11434 a_25019_n3588.t9 VSS 0.058887f
C11435 a_25019_n3588.t2 VSS 0.040077f
C11436 a_25019_n3588.n6 VSS 0.976326f
C11437 a_26060_n878.n0 VSS 11.128f
C11438 a_26060_n878.t0 VSS 0.295288f
C11439 a_26060_n878.t1 VSS 0.189924f
C11440 a_26060_n878.t3 VSS 0.247499f
C11441 a_26060_n878.t2 VSS 0.297193f
C11442 a_26060_n878.n1 VSS 8.942089f
C11443 a_21996_n12996.t2 VSS 0.072606f
C11444 a_21996_n12996.n0 VSS 0.013063f
C11445 a_21996_n12996.t10 VSS 0.044893f
C11446 a_21996_n12996.t8 VSS 0.03653f
C11447 a_21996_n12996.n1 VSS 0.076826f
C11448 a_21996_n12996.t4 VSS 0.03653f
C11449 a_21996_n12996.t12 VSS 0.044893f
C11450 a_21996_n12996.n2 VSS 0.117861f
C11451 a_21996_n12996.t6 VSS 0.044893f
C11452 a_21996_n12996.t7 VSS 0.03653f
C11453 a_21996_n12996.n3 VSS 0.092162f
C11454 a_21996_n12996.n4 VSS 0.690111f
C11455 a_21996_n12996.t5 VSS 0.044893f
C11456 a_21996_n12996.t9 VSS 0.03653f
C11457 a_21996_n12996.n5 VSS 0.076701f
C11458 a_21996_n12996.n6 VSS 0.585989f
C11459 a_21996_n12996.t11 VSS 0.044893f
C11460 a_21996_n12996.t3 VSS 0.03653f
C11461 a_21996_n12996.n7 VSS 0.076701f
C11462 a_21996_n12996.n8 VSS 0.569722f
C11463 a_21996_n12996.n9 VSS 1.20937f
C11464 a_21996_n12996.n10 VSS 0.70044f
C11465 a_28009_n1192.t1 VSS 7.60413f
C11466 a_28009_n1192.t2 VSS 0.154989f
C11467 a_28009_n1192.t3 VSS 0.199256f
C11468 a_28009_n1192.n0 VSS 5.7136f
C11469 a_28009_n1192.t0 VSS 0.128019f
C11470 a_23564_n14564.t1 VSS 1.31517f
C11471 a_23564_n14564.n0 VSS 0.111464f
C11472 a_23564_n14564.t0 VSS 0.03794f
C11473 a_23564_n14564.t5 VSS 0.060065f
C11474 a_23564_n14564.t9 VSS 0.055417f
C11475 a_23564_n14564.n1 VSS 0.09184f
C11476 a_23564_n14564.t3 VSS 0.060065f
C11477 a_23564_n14564.t4 VSS 0.062295f
C11478 a_23564_n14564.t8 VSS 0.052571f
C11479 a_23564_n14564.n2 VSS 0.09739f
C11480 a_23564_n14564.t6 VSS 0.052571f
C11481 a_23564_n14564.t7 VSS 0.060065f
C11482 a_23564_n14564.t2 VSS 0.055417f
C11483 a_23564_n14564.n3 VSS 1.18773f
C11484 a_23564_1116.t1 VSS 17.1575f
C11485 a_23564_1116.n0 VSS 0.654446f
C11486 a_23564_1116.t0 VSS 0.22563f
C11487 a_23564_1116.t9 VSS 0.352662f
C11488 a_23564_1116.t5 VSS 0.325377f
C11489 a_23564_1116.n1 VSS 0.539227f
C11490 a_23564_1116.t7 VSS 0.352662f
C11491 a_23564_1116.t8 VSS 0.36576f
C11492 a_23564_1116.t4 VSS 0.308662f
C11493 a_23564_1116.n2 VSS 0.571815f
C11494 a_23564_1116.t3 VSS 0.308662f
C11495 a_23564_1116.t2 VSS 0.352662f
C11496 a_23564_1116.t6 VSS 0.325377f
C11497 a_23564_1116.n3 VSS 15.159499f
C11498 a_22724_860.t1 VSS 0.421531f
C11499 a_22724_860.t0 VSS 0.038068f
C11500 a_22724_860.t6 VSS 0.175684f
C11501 a_22724_860.t4 VSS 0.231525f
C11502 a_22724_860.t3 VSS 0.13409f
C11503 a_22724_860.t2 VSS 0.450407f
C11504 a_22724_860.t5 VSS 0.539579f
C11505 a_22724_860.t7 VSS 0.293265f
C11506 a_22724_860.n0 VSS 0.115851f
C11507 a_21804_n2273.n0 VSS 1.28527f
C11508 a_21804_n2273.t1 VSS 0.824773f
C11509 a_21804_n2273.t0 VSS 0.042729f
C11510 a_21804_n2273.t11 VSS 0.028877f
C11511 a_21804_n2273.t13 VSS 0.031598f
C11512 a_21804_n2273.n1 VSS 0.465465f
C11513 a_21804_n2273.t12 VSS 0.036313f
C11514 a_21804_n2273.t3 VSS 0.068934f
C11515 a_21804_n2273.n2 VSS 0.195196f
C11516 a_21804_n2273.t9 VSS 0.028877f
C11517 a_21804_n2273.t8 VSS 0.031598f
C11518 a_21804_n2273.t2 VSS 0.068934f
C11519 a_21804_n2273.t6 VSS 0.036313f
C11520 a_21804_n2273.n3 VSS 0.073571f
C11521 a_21804_n2273.t4 VSS 0.032207f
C11522 a_21804_n2273.t5 VSS 0.028868f
C11523 a_21804_n2273.n4 VSS 0.34284f
C11524 a_21804_n2273.n5 VSS 0.806337f
C11525 a_21804_n2273.t7 VSS 0.062955f
C11526 a_21804_n2273.t10 VSS 0.065907f
C11527 a_21804_n2273.n6 VSS 0.077009f
C11528 a_21804_n2273.n7 VSS 1.1384f
C11529 a_21804_n2273.n8 VSS 1.73963f
C11530 a_21804_n2273.n9 VSS 2.2874f
C11531 a_24716_n5156.t0 VSS 0.023827f
C11532 a_24716_n5156.t5 VSS 0.038401f
C11533 a_24716_n5156.t7 VSS 0.018973f
C11534 a_24716_n5156.n0 VSS 0.152502f
C11535 a_24716_n5156.t4 VSS 0.043329f
C11536 a_24716_n5156.t3 VSS 0.028441f
C11537 a_24716_n5156.n1 VSS 0.165077f
C11538 a_24716_n5156.t2 VSS 0.030528f
C11539 a_24716_n5156.t6 VSS 0.01944f
C11540 a_24716_n5156.n2 VSS 0.2742f
C11541 a_24716_n5156.n3 VSS 1.04712f
C11542 a_24716_n5156.n4 VSS 0.40622f
C11543 a_24716_n5156.n5 VSS 0.114126f
C11544 a_24716_n5156.t1 VSS 0.037812f
C11545 a_23564_n452.t1 VSS 8.4929f
C11546 a_23564_n452.n0 VSS 0.366766f
C11547 a_23564_n452.t0 VSS 0.070122f
C11548 a_23564_n452.t5 VSS 0.19764f
C11549 a_23564_n452.t7 VSS 0.182349f
C11550 a_23564_n452.n1 VSS 0.302195f
C11551 a_23564_n452.t3 VSS 0.19764f
C11552 a_23564_n452.t8 VSS 0.20498f
C11553 a_23564_n452.t6 VSS 0.172981f
C11554 a_23564_n452.n2 VSS 0.320458f
C11555 a_23564_n452.t4 VSS 0.172981f
C11556 a_23564_n452.t2 VSS 0.19764f
C11557 a_23564_n452.t9 VSS 0.182349f
C11558 a_23564_n452.n3 VSS 7.939f
C11559 a_21916_n6694.t0 VSS 0.103327f
C11560 a_21916_n6694.t1 VSS 0.168712f
C11561 a_21916_n6694.n0 VSS 0.32743f
C11562 a_21916_n6694.t9 VSS 0.087133f
C11563 a_21916_n6694.t21 VSS 0.100149f
C11564 a_21916_n6694.n1 VSS 0.493444f
C11565 a_21916_n6694.t2 VSS 0.1007f
C11566 a_21916_n6694.t19 VSS 0.075175f
C11567 a_21916_n6694.n2 VSS 0.482987f
C11568 a_21916_n6694.t18 VSS 0.098082f
C11569 a_21916_n6694.t17 VSS 0.104992f
C11570 a_21916_n6694.n3 VSS 0.209983f
C11571 a_21916_n6694.n4 VSS 1.92998f
C11572 a_21916_n6694.n5 VSS 1.63439f
C11573 a_21916_n6694.t11 VSS 0.072432f
C11574 a_21916_n6694.n6 VSS 0.068312f
C11575 a_21916_n6694.t15 VSS 0.094096f
C11576 a_21916_n6694.n7 VSS 0.107534f
C11577 a_21916_n6694.t8 VSS 0.094096f
C11578 a_21916_n6694.n8 VSS 0.107534f
C11579 a_21916_n6694.t13 VSS 0.072432f
C11580 a_21916_n6694.n9 VSS 0.066622f
C11581 a_21916_n6694.t10 VSS 0.072432f
C11582 a_21916_n6694.n10 VSS 0.068204f
C11583 a_21916_n6694.t16 VSS 0.094096f
C11584 a_21916_n6694.t4 VSS 0.094096f
C11585 a_21916_n6694.n11 VSS 0.107534f
C11586 a_21916_n6694.n12 VSS 0.107534f
C11587 a_21916_n6694.t12 VSS 0.072432f
C11588 a_21916_n6694.n13 VSS 0.066622f
C11589 a_21916_n6694.n14 VSS 0.813338f
C11590 a_21916_n6694.t14 VSS 0.102402f
C11591 a_21916_n6694.t5 VSS 0.092446f
C11592 a_21916_n6694.n15 VSS 0.135883f
C11593 a_21916_n6694.t3 VSS 0.077386f
C11594 a_21916_n6694.t7 VSS 0.113906f
C11595 a_21916_n6694.n16 VSS 0.130543f
C11596 a_21916_n6694.n17 VSS 0.152085f
C11597 a_21916_n6694.n18 VSS 0.933904f
C11598 a_21916_n6694.t6 VSS 0.090666f
C11599 a_21916_n6694.t20 VSS 0.104827f
C11600 a_21916_n6694.n19 VSS 0.375881f
C11601 a_21916_n6694.n20 VSS 1.65257f
C11602 a_21916_n6694.n21 VSS 0.441679f
C11603 a_n263_3472.n0 VSS 3.76518f
C11604 a_n263_3472.n1 VSS 0.076162f
C11605 a_n263_3472.t12 VSS 0.010498f
C11606 a_n263_3472.t11 VSS 0.010498f
C11607 a_n263_3472.t10 VSS 0.014536f
C11608 a_n263_3472.n2 VSS 0.025348f
C11609 a_n263_3472.t9 VSS 0.014536f
C11610 a_n263_3472.t8 VSS 0.010498f
C11611 a_n263_3472.n3 VSS 0.031615f
C11612 a_n263_3472.n4 VSS 0.014161f
C11613 a_n263_3472.n5 VSS 0.016971f
C11614 a_n263_3472.n6 VSS 0.014161f
C11615 a_n263_3472.n7 VSS 0.017027f
C11616 a_n263_3472.t14 VSS 0.010498f
C11617 a_n263_3472.t13 VSS 0.014536f
C11618 a_n263_3472.n8 VSS 0.025348f
C11619 a_n263_3472.t17 VSS 0.042686f
C11620 a_n263_3472.t18 VSS 0.041648f
C11621 a_n263_3472.n9 VSS 0.339446f
C11622 a_n263_3472.t16 VSS 0.048465f
C11623 a_n263_3472.n10 VSS 5.65985f
C11624 a_n263_3472.n11 VSS 0.025348f
C11625 a_n263_3472.t15 VSS 0.014536f
C11626 a_13501_n19850.n0 VSS 2.0189f
C11627 a_13501_n19850.n1 VSS 3.79312f
C11628 a_13501_n19850.t3 VSS 0.041646f
C11629 a_13501_n19850.t4 VSS 0.33153f
C11630 a_13501_n19850.t19 VSS 0.321965f
C11631 a_13501_n19850.t17 VSS 0.041646f
C11632 a_13501_n19850.t11 VSS 0.041646f
C11633 a_13501_n19850.n2 VSS 0.229216f
C11634 a_13501_n19850.t2 VSS 0.041646f
C11635 a_13501_n19850.t6 VSS 0.041646f
C11636 a_13501_n19850.n3 VSS 0.223712f
C11637 a_13501_n19850.t14 VSS 0.041646f
C11638 a_13501_n19850.t18 VSS 0.041646f
C11639 a_13501_n19850.n4 VSS 0.228449f
C11640 a_13501_n19850.t5 VSS 0.33124f
C11641 a_13501_n19850.t10 VSS 0.325425f
C11642 a_13501_n19850.t8 VSS 0.041646f
C11643 a_13501_n19850.t1 VSS 0.041646f
C11644 a_13501_n19850.n5 VSS 0.22387f
C11645 a_13501_n19850.t13 VSS 0.041646f
C11646 a_13501_n19850.t16 VSS 0.041646f
C11647 a_13501_n19850.n6 VSS 0.228065f
C11648 a_13501_n19850.t12 VSS 0.041646f
C11649 a_13501_n19850.t15 VSS 0.041646f
C11650 a_13501_n19850.n7 VSS 0.227874f
C11651 a_13501_n19850.t7 VSS 0.041646f
C11652 a_13501_n19850.t0 VSS 0.041646f
C11653 a_13501_n19850.n8 VSS 0.22515f
C11654 a_13501_n19850.n9 VSS 0.22515f
C11655 a_13501_n19850.t9 VSS 0.041646f
C11656 a_41392_1944.n0 VSS 0.400016f
C11657 a_41392_1944.t4 VSS 0.020507f
C11658 a_41392_1944.t6 VSS 0.028394f
C11659 a_41392_1944.t5 VSS 0.020507f
C11660 a_41392_1944.n1 VSS 0.049378f
C11661 a_41392_1944.t2 VSS 0.013783f
C11662 a_41392_1944.t1 VSS 0.013783f
C11663 a_41392_1944.n2 VSS 0.027645f
C11664 a_41392_1944.t3 VSS 0.013783f
C11665 a_41392_1944.t0 VSS 0.013783f
C11666 a_41392_1944.n3 VSS 0.033293f
C11667 a_41392_1944.t18 VSS 0.057602f
C11668 a_41392_1944.t10 VSS 0.06058f
C11669 a_41392_1944.n4 VSS 0.094008f
C11670 a_41392_1944.t21 VSS 0.057602f
C11671 a_41392_1944.t13 VSS 0.06058f
C11672 a_41392_1944.n5 VSS -0.036634f
C11673 a_41392_1944.t17 VSS 0.057602f
C11674 a_41392_1944.t9 VSS 0.06058f
C11675 a_41392_1944.n6 VSS 0.10611f
C11676 a_41392_1944.t23 VSS 0.057602f
C11677 a_41392_1944.t15 VSS 0.06058f
C11678 a_41392_1944.n7 VSS 0.10611f
C11679 a_41392_1944.t20 VSS 0.057602f
C11680 a_41392_1944.t12 VSS 0.06058f
C11681 a_41392_1944.n8 VSS 0.10611f
C11682 a_41392_1944.t16 VSS 0.057602f
C11683 a_41392_1944.t8 VSS 0.06058f
C11684 a_41392_1944.n9 VSS 0.10611f
C11685 a_41392_1944.t22 VSS 0.057602f
C11686 a_41392_1944.t14 VSS 0.06058f
C11687 a_41392_1944.n10 VSS 0.094008f
C11688 a_41392_1944.t19 VSS 0.057602f
C11689 a_41392_1944.t11 VSS 0.06058f
C11690 a_41392_1944.n11 VSS 0.152616f
C11691 a_41392_1944.n12 VSS 0.06284f
C11692 a_41392_1944.t7 VSS 0.028394f
C11693 a_29532_n4372.n0 VSS 0.560575f
C11694 a_29532_n4372.t3 VSS 0.054093f
C11695 a_29532_n4372.t0 VSS 0.063713f
C11696 a_29532_n4372.t2 VSS 0.059223f
C11697 a_29532_n4372.t1 VSS 0.059223f
C11698 a_29532_n4372.t5 VSS 0.054225f
C11699 a_29532_n4372.t7 VSS 0.051511f
C11700 a_29532_n4372.n1 VSS 0.348293f
C11701 a_29532_n4372.t8 VSS 0.055891f
C11702 a_29532_n4372.t9 VSS 0.046106f
C11703 a_29532_n4372.n2 VSS 0.070924f
C11704 a_29532_n4372.t6 VSS 0.070978f
C11705 a_29532_n4372.t4 VSS 0.031941f
C11706 a_29532_n4372.n3 VSS 0.088952f
C11707 a_29532_n4372.n4 VSS 0.235845f
C11708 a_29532_n4372.n5 VSS 0.948506f
C11709 OUT[0].t6 VSS 0.015262f
C11710 OUT[0].t3 VSS 0.015262f
C11711 OUT[0].n0 VSS 0.03063f
C11712 OUT[0].t2 VSS 0.015262f
C11713 OUT[0].t0 VSS 0.015262f
C11714 OUT[0].n1 VSS 0.03063f
C11715 OUT[0].t1 VSS 0.015262f
C11716 OUT[0].t5 VSS 0.015262f
C11717 OUT[0].n2 VSS 0.036706f
C11718 OUT[0].n3 VSS 0.167641f
C11719 OUT[0].t14 VSS 0.031441f
C11720 OUT[0].t11 VSS 0.022708f
C11721 OUT[0].n4 VSS 0.054828f
C11722 OUT[0].t15 VSS 0.022708f
C11723 OUT[0].t12 VSS 0.031441f
C11724 OUT[0].n5 VSS 0.068381f
C11725 OUT[0].n6 VSS 0.172031f
C11726 OUT[0].t10 VSS 0.031441f
C11727 OUT[0].t8 VSS 0.022708f
C11728 OUT[0].n7 VSS 0.054828f
C11729 OUT[0].t9 VSS 0.031441f
C11730 OUT[0].t13 VSS 0.022708f
C11731 OUT[0].n8 VSS 0.069357f
C11732 OUT[0].n9 VSS 0.175408f
C11733 OUT[0].n10 VSS 0.134813f
C11734 OUT[0].n11 VSS 0.134813f
C11735 OUT[0].n12 VSS 0.096161f
C11736 OUT[0].t7 VSS 0.015262f
C11737 OUT[0].t4 VSS 0.015262f
C11738 OUT[0].n13 VSS 0.030525f
C11739 OUT[0].n14 VSS 0.329051f
C11740 a_29408_1944.n0 VSS 0.383348f
C11741 a_29408_1944.t5 VSS 0.027211f
C11742 a_29408_1944.t4 VSS 0.027211f
C11743 a_29408_1944.t6 VSS 0.019652f
C11744 a_29408_1944.n1 VSS 0.047321f
C11745 a_29408_1944.t0 VSS 0.013209f
C11746 a_29408_1944.t2 VSS 0.013209f
C11747 a_29408_1944.n2 VSS 0.026494f
C11748 a_29408_1944.t1 VSS 0.013209f
C11749 a_29408_1944.t3 VSS 0.013209f
C11750 a_29408_1944.n3 VSS 0.031906f
C11751 a_29408_1944.t14 VSS 0.055202f
C11752 a_29408_1944.t22 VSS 0.058056f
C11753 a_29408_1944.n4 VSS 0.090091f
C11754 a_29408_1944.t10 VSS 0.055202f
C11755 a_29408_1944.t18 VSS 0.058056f
C11756 a_29408_1944.n5 VSS -0.035108f
C11757 a_29408_1944.t13 VSS 0.055202f
C11758 a_29408_1944.t21 VSS 0.058056f
C11759 a_29408_1944.n6 VSS 0.101689f
C11760 a_29408_1944.t15 VSS 0.055202f
C11761 a_29408_1944.t23 VSS 0.058056f
C11762 a_29408_1944.n7 VSS 0.101689f
C11763 a_29408_1944.t9 VSS 0.055202f
C11764 a_29408_1944.t17 VSS 0.058056f
C11765 a_29408_1944.n8 VSS 0.101689f
C11766 a_29408_1944.t12 VSS 0.055202f
C11767 a_29408_1944.t20 VSS 0.058056f
C11768 a_29408_1944.n9 VSS 0.101689f
C11769 a_29408_1944.t11 VSS 0.055202f
C11770 a_29408_1944.t19 VSS 0.058056f
C11771 a_29408_1944.n10 VSS 0.090091f
C11772 a_29408_1944.t8 VSS 0.055202f
C11773 a_29408_1944.t16 VSS 0.058056f
C11774 a_29408_1944.n11 VSS 0.146257f
C11775 a_29408_1944.n12 VSS 0.060222f
C11776 a_29408_1944.t7 VSS 0.019652f
C11777 a_22444_2253.n0 VSS 0.400114f
C11778 a_22444_2253.t6 VSS 0.028394f
C11779 a_22444_2253.t4 VSS 0.020507f
C11780 a_22444_2253.t5 VSS 0.028394f
C11781 a_22444_2253.n1 VSS 0.049378f
C11782 a_22444_2253.t0 VSS 0.013783f
C11783 a_22444_2253.t2 VSS 0.013783f
C11784 a_22444_2253.n2 VSS 0.027645f
C11785 a_22444_2253.t3 VSS 0.013783f
C11786 a_22444_2253.t1 VSS 0.013783f
C11787 a_22444_2253.n3 VSS 0.033293f
C11788 a_22444_2253.t22 VSS 0.057602f
C11789 a_22444_2253.t20 VSS 0.06058f
C11790 a_22444_2253.n4 VSS 0.094008f
C11791 a_22444_2253.t14 VSS 0.057602f
C11792 a_22444_2253.t11 VSS 0.06058f
C11793 a_22444_2253.n5 VSS 0.094008f
C11794 a_22444_2253.t10 VSS 0.057602f
C11795 a_22444_2253.t9 VSS 0.06058f
C11796 a_22444_2253.n6 VSS -0.036634f
C11797 a_22444_2253.t17 VSS 0.057602f
C11798 a_22444_2253.t8 VSS 0.06058f
C11799 a_22444_2253.n7 VSS 0.10611f
C11800 a_22444_2253.t16 VSS 0.057602f
C11801 a_22444_2253.t13 VSS 0.06058f
C11802 a_22444_2253.n8 VSS 0.10611f
C11803 a_22444_2253.t21 VSS 0.057602f
C11804 a_22444_2253.t19 VSS 0.06058f
C11805 a_22444_2253.n9 VSS 0.10611f
C11806 a_22444_2253.t18 VSS 0.057602f
C11807 a_22444_2253.t15 VSS 0.06058f
C11808 a_22444_2253.n10 VSS 0.10611f
C11809 a_22444_2253.t12 VSS 0.057602f
C11810 a_22444_2253.t23 VSS 0.06058f
C11811 a_22444_2253.n11 VSS 0.152517f
C11812 a_22444_2253.n12 VSS 0.06284f
C11813 a_22444_2253.t7 VSS 0.020507f
C11814 a_24236_2258.t1 VSS 2.45863f
C11815 a_24236_2258.n0 VSS 0.089899f
C11816 a_24236_2258.t0 VSS 0.017188f
C11817 a_24236_2258.t3 VSS 0.044696f
C11818 a_24236_2258.t2 VSS 0.048444f
C11819 a_24236_2258.n1 VSS 0.074072f
C11820 a_24236_2258.t6 VSS 0.0424f
C11821 a_24236_2258.t5 VSS 0.050243f
C11822 a_24236_2258.n2 VSS 0.078548f
C11823 a_24236_2258.t9 VSS 0.0424f
C11824 a_24236_2258.t8 VSS 0.048444f
C11825 a_24236_2258.t7 VSS 0.044696f
C11826 a_24236_2258.t4 VSS 0.048444f
C11827 a_24236_2258.n3 VSS 2.2119f
C11828 a_1955_4292.t3 VSS 0.040666f
C11829 a_1955_4292.t2 VSS 0.053922f
C11830 a_1955_4292.t4 VSS 0.046744f
C11831 a_1955_4292.n0 VSS 0.539245f
C11832 a_1955_4292.n1 VSS 0.999094f
C11833 a_1955_4292.t1 VSS 0.167423f
C11834 a_1955_4292.n2 VSS 1.52866f
C11835 a_1955_4292.t0 VSS 0.124245f
C11836 a_11023_n20230.n0 VSS 0.016619f
C11837 a_11023_n20230.n1 VSS 0.646071f
C11838 a_11023_n20230.n2 VSS 0.0574f
C11839 a_11023_n20230.n3 VSS 0.016723f
C11840 a_11023_n20230.n4 VSS 0.057191f
C11841 a_11023_n20230.n5 VSS 0.056982f
C11842 a_11023_n20230.n6 VSS 0.056773f
C11843 a_11023_n20230.n7 VSS 0.318043f
C11844 a_11023_n20230.n8 VSS 0.318043f
C11845 a_11023_n20230.n9 VSS 0.318043f
C11846 a_11023_n20230.n10 VSS 0.440197f
C11847 a_11023_n20230.n11 VSS 0.107951f
C11848 a_11023_n20230.n12 VSS 0.052801f
C11849 a_11023_n20230.n13 VSS 0.022159f
C11850 a_11023_n20230.n14 VSS 0.052592f
C11851 a_11023_n20230.n15 VSS 0.022159f
C11852 a_11023_n20230.n16 VSS 0.052383f
C11853 a_11023_n20230.n17 VSS 0.052174f
C11854 a_11023_n20230.t12 VSS 0.038046f
C11855 a_11023_n20230.t17 VSS 0.038046f
C11856 a_11023_n20230.t11 VSS 0.038046f
C11857 a_11023_n20230.n18 VSS 0.198238f
C11858 a_11023_n20230.t15 VSS 0.038046f
C11859 a_11023_n20230.t18 VSS 0.038046f
C11860 a_11023_n20230.n19 VSS 0.183088f
C11861 a_11023_n20230.n20 VSS 0.507916f
C11862 a_11023_n20230.t30 VSS 0.064777f
C11863 a_11023_n20230.n21 VSS 0.145665f
C11864 a_11023_n20230.t35 VSS 0.06465f
C11865 a_11023_n20230.n22 VSS 0.056431f
C11866 a_11023_n20230.t27 VSS 0.06465f
C11867 a_11023_n20230.n23 VSS 0.016723f
C11868 a_11023_n20230.n24 VSS 0.120365f
C11869 a_11023_n20230.n25 VSS 0.022159f
C11870 a_11023_n20230.n26 VSS 0.022159f
C11871 a_11023_n20230.t21 VSS 0.06465f
C11872 a_11023_n20230.t33 VSS 0.06465f
C11873 a_11023_n20230.t38 VSS 0.06465f
C11874 a_11023_n20230.t36 VSS 0.06465f
C11875 a_11023_n20230.t32 VSS 0.064506f
C11876 a_11023_n20230.t20 VSS 0.064403f
C11877 a_11023_n20230.t26 VSS 0.064403f
C11878 a_11023_n20230.t34 VSS 0.064403f
C11879 a_11023_n20230.t22 VSS 0.064403f
C11880 a_11023_n20230.t29 VSS 0.064403f
C11881 a_11023_n20230.t37 VSS 0.064403f
C11882 a_11023_n20230.t31 VSS 0.064403f
C11883 a_11023_n20230.t39 VSS 0.064403f
C11884 a_11023_n20230.t25 VSS 0.064403f
C11885 a_11023_n20230.n27 VSS 0.223528f
C11886 a_11023_n20230.t28 VSS 0.06465f
C11887 a_11023_n20230.n28 VSS 0.072599f
C11888 a_11023_n20230.n29 VSS 0.022159f
C11889 a_11023_n20230.n30 VSS 0.016723f
C11890 a_11023_n20230.t23 VSS 0.06465f
C11891 a_11023_n20230.n31 VSS 0.022159f
C11892 a_11023_n20230.n32 VSS 0.022159f
C11893 a_11023_n20230.n33 VSS 0.016723f
C11894 a_11023_n20230.t24 VSS 0.06465f
C11895 a_11023_n20230.t8 VSS 0.038046f
C11896 a_11023_n20230.t2 VSS 0.038046f
C11897 a_11023_n20230.n34 VSS 0.180651f
C11898 a_11023_n20230.t1 VSS 0.038046f
C11899 a_11023_n20230.t4 VSS 0.038046f
C11900 a_11023_n20230.n35 VSS 0.180651f
C11901 a_11023_n20230.t0 VSS 0.038046f
C11902 a_11023_n20230.t7 VSS 0.038046f
C11903 a_11023_n20230.n36 VSS 0.180651f
C11904 a_11023_n20230.t3 VSS 0.038046f
C11905 a_11023_n20230.t6 VSS 0.038046f
C11906 a_11023_n20230.n37 VSS 0.180651f
C11907 a_11023_n20230.t5 VSS 0.038046f
C11908 a_11023_n20230.t9 VSS 0.038046f
C11909 a_11023_n20230.n38 VSS 0.200645f
C11910 a_11023_n20230.n39 VSS 0.702578f
C11911 a_11023_n20230.n40 VSS 0.300774f
C11912 a_11023_n20230.n41 VSS 0.300774f
C11913 a_11023_n20230.n42 VSS 0.418266f
C11914 a_11023_n20230.n43 VSS 0.725258f
C11915 a_11023_n20230.t10 VSS 0.038046f
C11916 a_11023_n20230.t14 VSS 0.038046f
C11917 a_11023_n20230.n44 VSS 0.183088f
C11918 a_11023_n20230.n45 VSS 0.322395f
C11919 a_11023_n20230.t13 VSS 0.038046f
C11920 a_11023_n20230.t16 VSS 0.038046f
C11921 a_11023_n20230.n46 VSS 0.183088f
C11922 a_11023_n20230.n47 VSS 0.186332f
C11923 a_11023_n20230.n48 VSS 0.18633f
C11924 a_11023_n20230.n49 VSS 0.183091f
C11925 a_11023_n20230.t19 VSS 0.038046f
C11926 OUT[2].t1 VSS 0.013427f
C11927 OUT[2].t4 VSS 0.013427f
C11928 OUT[2].n0 VSS 0.026948f
C11929 OUT[2].t5 VSS 0.013427f
C11930 OUT[2].t7 VSS 0.013427f
C11931 OUT[2].n1 VSS 0.026948f
C11932 OUT[2].t3 VSS 0.013427f
C11933 OUT[2].t0 VSS 0.013427f
C11934 OUT[2].n2 VSS 0.032294f
C11935 OUT[2].n3 VSS 0.147487f
C11936 OUT[2].t10 VSS 0.027661f
C11937 OUT[2].t13 VSS 0.019978f
C11938 OUT[2].n4 VSS 0.048236f
C11939 OUT[2].t11 VSS 0.019978f
C11940 OUT[2].t15 VSS 0.027661f
C11941 OUT[2].n5 VSS 0.06016f
C11942 OUT[2].n6 VSS 0.151349f
C11943 OUT[2].t14 VSS 0.027661f
C11944 OUT[2].t8 VSS 0.019978f
C11945 OUT[2].n7 VSS 0.048236f
C11946 OUT[2].t12 VSS 0.027661f
C11947 OUT[2].t9 VSS 0.019978f
C11948 OUT[2].n8 VSS 0.061019f
C11949 OUT[2].n9 VSS 0.15432f
C11950 OUT[2].n10 VSS 0.118606f
C11951 OUT[2].n11 VSS 0.118606f
C11952 OUT[2].n12 VSS 0.084601f
C11953 OUT[2].t2 VSS 0.013427f
C11954 OUT[2].t6 VSS 0.013427f
C11955 OUT[2].n13 VSS 0.026855f
C11956 OUT[2].n14 VSS 0.415125f
C11957 a_37024_1944.n0 VSS 0.716695f
C11958 a_37024_1944.t4 VSS 0.036741f
C11959 a_37024_1944.t6 VSS 0.050872f
C11960 a_37024_1944.t5 VSS 0.036741f
C11961 a_37024_1944.n1 VSS 0.088469f
C11962 a_37024_1944.t1 VSS 0.024695f
C11963 a_37024_1944.t0 VSS 0.024695f
C11964 a_37024_1944.n2 VSS 0.049531f
C11965 a_37024_1944.t2 VSS 0.024695f
C11966 a_37024_1944.t3 VSS 0.024695f
C11967 a_37024_1944.n3 VSS 0.059649f
C11968 a_37024_1944.t19 VSS 0.103204f
C11969 a_37024_1944.t11 VSS 0.108539f
C11970 a_37024_1944.n4 VSS 0.168431f
C11971 a_37024_1944.t22 VSS 0.103204f
C11972 a_37024_1944.t14 VSS 0.108539f
C11973 a_37024_1944.n5 VSS -0.065636f
C11974 a_37024_1944.t17 VSS 0.103204f
C11975 a_37024_1944.t9 VSS 0.108539f
C11976 a_37024_1944.n6 VSS 0.190114f
C11977 a_37024_1944.t15 VSS 0.103204f
C11978 a_37024_1944.t23 VSS 0.108539f
C11979 a_37024_1944.n7 VSS 0.190114f
C11980 a_37024_1944.t21 VSS 0.103204f
C11981 a_37024_1944.t13 VSS 0.108539f
C11982 a_37024_1944.n8 VSS 0.190114f
C11983 a_37024_1944.t18 VSS 0.103204f
C11984 a_37024_1944.t10 VSS 0.108539f
C11985 a_37024_1944.n9 VSS 0.190114f
C11986 a_37024_1944.t16 VSS 0.103204f
C11987 a_37024_1944.t8 VSS 0.108539f
C11988 a_37024_1944.n10 VSS 0.168431f
C11989 a_37024_1944.t20 VSS 0.103204f
C11990 a_37024_1944.t12 VSS 0.108539f
C11991 a_37024_1944.n11 VSS 0.273436f
C11992 a_37024_1944.n12 VSS 0.112589f
C11993 a_37024_1944.t7 VSS 0.050872f
C11994 a_13623_n14874.n0 VSS 3.59854f
C11995 a_13623_n14874.n1 VSS 0.50879f
C11996 a_13623_n14874.n2 VSS 0.546795f
C11997 a_13623_n14874.n3 VSS 1.69261f
C11998 a_13623_n14874.n4 VSS 0.367787f
C11999 a_13623_n14874.t14 VSS 0.013423f
C12000 a_13623_n14874.t9 VSS 0.018586f
C12001 a_13623_n14874.t11 VSS 0.013423f
C12002 a_13623_n14874.n5 VSS 0.040422f
C12003 a_13623_n14874.t12 VSS 0.013423f
C12004 a_13623_n14874.t8 VSS 0.018586f
C12005 a_13623_n14874.n6 VSS 0.03241f
C12006 a_13623_n14874.t10 VSS 0.013423f
C12007 a_13623_n14874.t13 VSS 0.018586f
C12008 a_13623_n14874.n7 VSS 0.03354f
C12009 a_13623_n14874.t39 VSS 0.05215f
C12010 a_13623_n14874.t36 VSS 0.052349f
C12011 a_13623_n14874.t26 VSS 0.05215f
C12012 a_13623_n14874.t23 VSS 0.052349f
C12013 a_13623_n14874.t16 VSS 0.05215f
C12014 a_13623_n14874.t42 VSS 0.052349f
C12015 a_13623_n14874.t34 VSS 0.05215f
C12016 a_13623_n14874.t25 VSS 0.05215f
C12017 a_13623_n14874.t33 VSS 0.05215f
C12018 a_13623_n14874.t18 VSS 0.05215f
C12019 a_13623_n14874.t40 VSS 0.05215f
C12020 a_13623_n14874.t27 VSS 0.05215f
C12021 a_13623_n14874.t43 VSS 0.052447f
C12022 a_13623_n14874.t22 VSS 0.052339f
C12023 a_13623_n14874.t35 VSS 0.05215f
C12024 a_13623_n14874.t44 VSS 0.05215f
C12025 a_13623_n14874.t38 VSS 0.05215f
C12026 a_13623_n14874.t19 VSS 0.05215f
C12027 a_13623_n14874.t30 VSS 0.05215f
C12028 a_13623_n14874.t41 VSS 0.05215f
C12029 a_13623_n14874.t21 VSS 0.05215f
C12030 a_13623_n14874.t32 VSS 0.05215f
C12031 a_13623_n14874.t28 VSS 0.05215f
C12032 a_13623_n14874.t17 VSS 0.052175f
C12033 a_13623_n14874.t24 VSS 0.052349f
C12034 a_13623_n14874.t37 VSS 0.052349f
C12035 a_13623_n14874.t45 VSS 0.052349f
C12036 a_13623_n14874.t29 VSS 0.052349f
C12037 a_13623_n14874.t20 VSS 0.052349f
C12038 a_13623_n14874.t31 VSS 0.052349f
C12039 a_13623_n14874.n8 VSS 0.018106f
C12040 a_13623_n14874.n9 VSS 0.021698f
C12041 a_13623_n14874.n10 VSS 0.018106f
C12042 a_13623_n14874.n11 VSS 0.02177f
C12043 a_13623_n14874.n12 VSS 0.03241f
C12044 a_13623_n14874.t15 VSS 0.018586f
C12045 a_24348_n16087.t1 VSS 0.153931f
C12046 a_24348_n16087.t0 VSS 0.027278f
C12047 a_24348_n16087.t2 VSS 0.041773f
C12048 a_24348_n16087.t4 VSS 0.031185f
C12049 a_24348_n16087.n0 VSS 0.402771f
C12050 a_24348_n16087.t5 VSS 0.0396f
C12051 a_24348_n16087.t7 VSS 0.019566f
C12052 a_24348_n16087.n1 VSS 0.0967f
C12053 a_24348_n16087.n2 VSS 0.627838f
C12054 a_24348_n16087.t3 VSS 0.040425f
C12055 a_24348_n16087.t6 VSS 0.021295f
C12056 a_24348_n16087.n3 VSS 0.136361f
C12057 a_24348_n16087.n4 VSS 0.461276f
C12058 CLK.t12 VSS 0.033675f
C12059 CLK.t6 VSS 0.034379f
C12060 CLK.n0 VSS 0.100076f
C12061 CLK.t15 VSS 0.101757f
C12062 CLK.t8 VSS 0.067158f
C12063 CLK.t1 VSS 0.037339f
C12064 CLK.n1 VSS 0.18509f
C12065 CLK.t9 VSS 0.067158f
C12066 CLK.t3 VSS 0.037339f
C12067 CLK.n2 VSS 0.130731f
C12068 CLK.t4 VSS 0.097223f
C12069 CLK.t2 VSS 0.067158f
C12070 CLK.t10 VSS 0.037339f
C12071 CLK.n3 VSS 0.183843f
C12072 CLK.t5 VSS 0.067158f
C12073 CLK.t13 VSS 0.037339f
C12074 CLK.n4 VSS 0.130731f
C12075 CLK.t11 VSS 0.067158f
C12076 CLK.t14 VSS 0.037339f
C12077 CLK.n5 VSS 0.130731f
C12078 CLK.t7 VSS 0.067158f
C12079 CLK.t0 VSS 0.037339f
C12080 CLK.n6 VSS 0.60105f
C12081 CLK.n7 VSS 2.01902f
C12082 a_13623_n12196.n0 VSS 3.63501f
C12083 a_13623_n12196.n1 VSS 0.543853f
C12084 a_13623_n12196.n2 VSS 0.584478f
C12085 a_13623_n12196.n3 VSS 1.52122f
C12086 a_13623_n12196.n4 VSS 0.393134f
C12087 a_13623_n12196.t14 VSS 0.014348f
C12088 a_13623_n12196.t9 VSS 0.019867f
C12089 a_13623_n12196.t11 VSS 0.014348f
C12090 a_13623_n12196.n5 VSS 0.043208f
C12091 a_13623_n12196.t12 VSS 0.014348f
C12092 a_13623_n12196.t8 VSS 0.019867f
C12093 a_13623_n12196.n6 VSS 0.034644f
C12094 a_13623_n12196.t10 VSS 0.014348f
C12095 a_13623_n12196.t13 VSS 0.019867f
C12096 a_13623_n12196.n7 VSS 0.035852f
C12097 a_13623_n12196.t40 VSS 0.055744f
C12098 a_13623_n12196.t43 VSS 0.055957f
C12099 a_13623_n12196.t26 VSS 0.055744f
C12100 a_13623_n12196.t31 VSS 0.055957f
C12101 a_13623_n12196.t16 VSS 0.055744f
C12102 a_13623_n12196.t20 VSS 0.055957f
C12103 a_13623_n12196.t35 VSS 0.055744f
C12104 a_13623_n12196.t25 VSS 0.055744f
C12105 a_13623_n12196.t34 VSS 0.055744f
C12106 a_13623_n12196.t18 VSS 0.055744f
C12107 a_13623_n12196.t41 VSS 0.055744f
C12108 a_13623_n12196.t27 VSS 0.055744f
C12109 a_13623_n12196.t21 VSS 0.056062f
C12110 a_13623_n12196.t23 VSS 0.055946f
C12111 a_13623_n12196.t36 VSS 0.055744f
C12112 a_13623_n12196.t45 VSS 0.055744f
C12113 a_13623_n12196.t38 VSS 0.055744f
C12114 a_13623_n12196.t19 VSS 0.055744f
C12115 a_13623_n12196.t30 VSS 0.055744f
C12116 a_13623_n12196.t42 VSS 0.055744f
C12117 a_13623_n12196.t22 VSS 0.055744f
C12118 a_13623_n12196.t33 VSS 0.055744f
C12119 a_13623_n12196.t28 VSS 0.055744f
C12120 a_13623_n12196.t17 VSS 0.055771f
C12121 a_13623_n12196.t32 VSS 0.055957f
C12122 a_13623_n12196.t44 VSS 0.055957f
C12123 a_13623_n12196.t24 VSS 0.055957f
C12124 a_13623_n12196.t37 VSS 0.055957f
C12125 a_13623_n12196.t29 VSS 0.055957f
C12126 a_13623_n12196.t39 VSS 0.055957f
C12127 a_13623_n12196.n8 VSS 0.019354f
C12128 a_13623_n12196.n9 VSS 0.023194f
C12129 a_13623_n12196.n10 VSS 0.019354f
C12130 a_13623_n12196.n11 VSS 0.02327f
C12131 a_13623_n12196.n12 VSS 0.034644f
C12132 a_13623_n12196.t15 VSS 0.019867f
C12133 a_21772_n14564.n0 VSS 0.61362f
C12134 a_21772_n14564.t3 VSS 0.055212f
C12135 a_21772_n14564.t0 VSS 0.060859f
C12136 a_21772_n14564.t1 VSS 0.067887f
C12137 a_21772_n14564.t2 VSS 0.081141f
C12138 a_21772_n14564.t14 VSS 0.06058f
C12139 a_21772_n14564.t4 VSS 0.057602f
C12140 a_21772_n14564.n1 VSS 0.094008f
C12141 a_21772_n14564.t8 VSS 0.06058f
C12142 a_21772_n14564.t17 VSS 0.057602f
C12143 a_21772_n14564.n2 VSS 0.094008f
C12144 a_21772_n14564.t12 VSS 0.06058f
C12145 a_21772_n14564.t10 VSS 0.057602f
C12146 a_21772_n14564.n3 VSS -0.036634f
C12147 a_21772_n14564.t15 VSS 0.06058f
C12148 a_21772_n14564.t5 VSS 0.057602f
C12149 a_21772_n14564.n4 VSS 0.106111f
C12150 a_21772_n14564.t9 VSS 0.06058f
C12151 a_21772_n14564.t18 VSS 0.057602f
C12152 a_21772_n14564.n5 VSS 0.106111f
C12153 a_21772_n14564.t6 VSS 0.06058f
C12154 a_21772_n14564.t13 VSS 0.057602f
C12155 a_21772_n14564.n6 VSS 0.106111f
C12156 a_21772_n14564.t7 VSS 0.06058f
C12157 a_21772_n14564.t16 VSS 0.057602f
C12158 a_21772_n14564.n7 VSS 0.106111f
C12159 a_21772_n14564.t11 VSS 0.06058f
C12160 a_21772_n14564.t19 VSS 0.057602f
C12161 a_29744_n15604.n0 VSS 0.448816f
C12162 a_29744_n15604.t4 VSS 0.023188f
C12163 a_29744_n15604.t1 VSS 0.020552f
C12164 a_29744_n15604.n1 VSS 0.024427f
C12165 a_29744_n15604.t21 VSS 0.073413f
C12166 a_29744_n15604.t14 VSS 0.044539f
C12167 a_29744_n15604.n2 VSS 0.106957f
C12168 a_29744_n15604.t20 VSS 0.073413f
C12169 a_29744_n15604.t10 VSS 0.044539f
C12170 a_29744_n15604.n3 VSS -0.028686f
C12171 a_29744_n15604.t16 VSS 0.073413f
C12172 a_29744_n15604.t8 VSS 0.044539f
C12173 a_29744_n15604.n4 VSS 0.121662f
C12174 a_29744_n15604.t22 VSS 0.073413f
C12175 a_29744_n15604.t13 VSS 0.044539f
C12176 a_29744_n15604.n5 VSS 0.121662f
C12177 a_29744_n15604.t18 VSS 0.073413f
C12178 a_29744_n15604.t12 VSS 0.044539f
C12179 a_29744_n15604.n6 VSS 0.121662f
C12180 a_29744_n15604.t7 VSS 0.073413f
C12181 a_29744_n15604.t15 VSS 0.044539f
C12182 a_29744_n15604.n7 VSS 0.118692f
C12183 a_29744_n15604.t19 VSS 0.073413f
C12184 a_29744_n15604.t9 VSS 0.044539f
C12185 a_29744_n15604.n8 VSS 0.106957f
C12186 a_29744_n15604.t17 VSS 0.073413f
C12187 a_29744_n15604.t11 VSS 0.044539f
C12188 a_29744_n15604.n9 VSS 0.109926f
C12189 a_29744_n15604.n10 VSS 0.071373f
C12190 a_29744_n15604.t3 VSS 0.023188f
C12191 a_29744_n15604.t5 VSS 0.023188f
C12192 a_29744_n15604.n11 VSS 0.056236f
C12193 a_29744_n15604.n12 VSS 0.046856f
C12194 a_29744_n15604.t6 VSS 0.023188f
C12195 a_21772_n17700.n0 VSS 0.38344f
C12196 a_21772_n17700.t6 VSS 0.027211f
C12197 a_21772_n17700.t5 VSS 0.019652f
C12198 a_21772_n17700.t4 VSS 0.027211f
C12199 a_21772_n17700.n1 VSS 0.060222f
C12200 a_21772_n17700.t2 VSS 0.013209f
C12201 a_21772_n17700.t1 VSS 0.013209f
C12202 a_21772_n17700.n2 VSS 0.026494f
C12203 a_21772_n17700.t0 VSS 0.013209f
C12204 a_21772_n17700.t3 VSS 0.013209f
C12205 a_21772_n17700.n3 VSS 0.031906f
C12206 a_21772_n17700.t18 VSS 0.058056f
C12207 a_21772_n17700.t8 VSS 0.055202f
C12208 a_21772_n17700.n4 VSS 0.090091f
C12209 a_21772_n17700.t12 VSS 0.058056f
C12210 a_21772_n17700.t21 VSS 0.055202f
C12211 a_21772_n17700.n5 VSS 0.090091f
C12212 a_21772_n17700.t16 VSS 0.058056f
C12213 a_21772_n17700.t14 VSS 0.055202f
C12214 a_21772_n17700.n6 VSS -0.035108f
C12215 a_21772_n17700.t19 VSS 0.058056f
C12216 a_21772_n17700.t9 VSS 0.055202f
C12217 a_21772_n17700.n7 VSS 0.101689f
C12218 a_21772_n17700.t13 VSS 0.058056f
C12219 a_21772_n17700.t22 VSS 0.055202f
C12220 a_21772_n17700.n8 VSS 0.101689f
C12221 a_21772_n17700.t10 VSS 0.058056f
C12222 a_21772_n17700.t17 VSS 0.055202f
C12223 a_21772_n17700.n9 VSS 0.101689f
C12224 a_21772_n17700.t11 VSS 0.058056f
C12225 a_21772_n17700.t20 VSS 0.055202f
C12226 a_21772_n17700.n10 VSS 0.101689f
C12227 a_21772_n17700.t15 VSS 0.058056f
C12228 a_21772_n17700.t23 VSS 0.055202f
C12229 a_21772_n17700.n11 VSS 0.146163f
C12230 a_21772_n17700.n12 VSS 0.047321f
C12231 a_21772_n17700.t7 VSS 0.019652f
C12232 a_30192_n15304.n0 VSS 0.466769f
C12233 a_30192_n15304.t4 VSS 0.024116f
C12234 a_30192_n15304.t5 VSS 0.024116f
C12235 a_30192_n15304.t3 VSS 0.024116f
C12236 a_30192_n15304.n1 VSS 0.04873f
C12237 a_30192_n15304.t2 VSS 0.021374f
C12238 a_30192_n15304.n2 VSS 0.025404f
C12239 a_30192_n15304.t18 VSS 0.04632f
C12240 a_30192_n15304.t8 VSS 0.076349f
C12241 a_30192_n15304.n3 VSS 0.111235f
C12242 a_30192_n15304.t16 VSS 0.04632f
C12243 a_30192_n15304.t10 VSS 0.076349f
C12244 a_30192_n15304.n4 VSS -0.029833f
C12245 a_30192_n15304.t21 VSS 0.04632f
C12246 a_30192_n15304.t11 VSS 0.076349f
C12247 a_30192_n15304.n5 VSS 0.126528f
C12248 a_30192_n15304.t15 VSS 0.04632f
C12249 a_30192_n15304.t9 VSS 0.076349f
C12250 a_30192_n15304.n6 VSS 0.126528f
C12251 a_30192_n15304.t14 VSS 0.04632f
C12252 a_30192_n15304.t20 VSS 0.076349f
C12253 a_30192_n15304.n7 VSS 0.126528f
C12254 a_30192_n15304.t19 VSS 0.04632f
C12255 a_30192_n15304.t12 VSS 0.076349f
C12256 a_30192_n15304.n8 VSS 0.12344f
C12257 a_30192_n15304.t22 VSS 0.04632f
C12258 a_30192_n15304.t13 VSS 0.076349f
C12259 a_30192_n15304.n9 VSS 0.111235f
C12260 a_30192_n15304.t17 VSS 0.04632f
C12261 a_30192_n15304.t7 VSS 0.076349f
C12262 a_30192_n15304.n10 VSS 0.114323f
C12263 a_30192_n15304.n11 VSS 0.074228f
C12264 a_30192_n15304.n12 VSS 0.058485f
C12265 a_30192_n15304.t6 VSS 0.024116f
C12266 a_11087_n20850.t31 VSS 6.81261f
C12267 a_11087_n20850.n0 VSS 0.19977f
C12268 a_11087_n20850.t37 VSS 2.71674f
C12269 a_11087_n20850.t32 VSS 5.72663f
C12270 a_11087_n20850.n1 VSS 1.0318f
C12271 a_11087_n20850.n2 VSS 0.358828f
C12272 a_11087_n20850.n3 VSS 1.88088f
C12273 a_11087_n20850.t30 VSS 3.40287f
C12274 a_11087_n20850.t41 VSS 2.14625f
C12275 a_11087_n20850.t36 VSS 2.21462f
C12276 a_11087_n20850.n4 VSS 0.355857f
C12277 a_11087_n20850.t38 VSS 3.40287f
C12278 a_11087_n20850.n5 VSS 0.020592f
C12279 a_11087_n20850.n6 VSS 0.026159f
C12280 a_11087_n20850.t34 VSS 2.64629f
C12281 a_11087_n20850.t33 VSS 2.73828f
C12282 a_11087_n20850.n7 VSS 0.020592f
C12283 a_11087_n20850.t35 VSS 1.27255f
C12284 a_11087_n20850.n8 VSS 1.08376f
C12285 a_11087_n20850.n9 VSS 0.020592f
C12286 a_11087_n20850.n10 VSS 0.032917f
C12287 a_11087_n20850.n11 VSS 0.029682f
C12288 a_11087_n20850.n12 VSS 0.022789f
C12289 a_11087_n20850.n13 VSS 0.012014f
C12290 a_11087_n20850.n14 VSS 0.032917f
C12291 a_11087_n20850.n15 VSS 0.49293f
C12292 a_11087_n20850.n16 VSS 0.020592f
C12293 a_11087_n20850.n17 VSS 0.014873f
C12294 a_11087_n20850.n18 VSS 0.012014f
C12295 a_11087_n20850.n19 VSS 0.012014f
C12296 a_11087_n20850.n20 VSS 0.012014f
C12297 a_11087_n20850.n21 VSS 0.06786f
C12298 a_11087_n20850.t7 VSS 0.053938f
C12299 a_11087_n20850.t10 VSS 0.055695f
C12300 a_11087_n20850.t29 VSS 0.054972f
C12301 a_11087_n20850.t21 VSS 0.053651f
C12302 a_11087_n20850.n22 VSS 0.153005f
C12303 a_11087_n20850.t28 VSS 0.053398f
C12304 a_11087_n20850.n23 VSS 0.05229f
C12305 a_11087_n20850.t25 VSS 0.053879f
C12306 a_11087_n20850.n24 VSS 0.052776f
C12307 a_11087_n20850.t26 VSS 0.053398f
C12308 a_11087_n20850.n25 VSS 0.092043f
C12309 a_11087_n20850.t40 VSS 2.44411f
C12310 a_11087_n20850.n26 VSS 0.357708f
C12311 a_11087_n20850.t39 VSS 2.39761f
C12312 a_11087_n20850.n27 VSS 0.032986f
C12313 a_11087_n20850.n28 VSS 0.056432f
C12314 a_11087_n20850.n29 VSS 0.043115f
C12315 a_11087_n20850.n30 VSS 0.043046f
C12316 a_11087_n20850.n31 VSS 0.032986f
C12317 a_11087_n20850.n32 VSS 0.015422f
C12318 a_11087_n20850.n33 VSS 0.015965f
C12319 a_11087_n20850.n34 VSS 0.023111f
C12320 a_11087_n20850.n35 VSS 0.041364f
C12321 a_11087_n20850.n36 VSS 0.015549f
C12322 a_11087_n20850.n37 VSS 0.138726f
C12323 a_11087_n20850.n38 VSS 0.358568f
C12324 a_11087_n20850.n39 VSS 0.830499f
C12325 a_11087_n20850.t0 VSS 0.054659f
C12326 a_11087_n20850.n40 VSS 0.179277f
C12327 a_11087_n20850.t14 VSS 0.054659f
C12328 a_11087_n20850.n41 VSS 0.045324f
C12329 a_11087_n20850.t9 VSS 0.053884f
C12330 a_11087_n20850.n42 VSS 0.044923f
C12331 a_11087_n20850.t11 VSS 0.053884f
C12332 a_11087_n20850.n43 VSS 0.045156f
C12333 a_11087_n20850.t5 VSS 0.053884f
C12334 a_11087_n20850.n44 VSS 0.06122f
C12335 a_11087_n20850.n45 VSS 0.1896f
C12336 a_11087_n20850.t16 VSS 0.054542f
C12337 a_11087_n20850.n46 VSS 0.121737f
C12338 a_11087_n20850.t18 VSS 0.054369f
C12339 a_11087_n20850.n47 VSS 0.044802f
C12340 a_11087_n20850.t13 VSS 0.054542f
C12341 a_11087_n20850.n48 VSS 0.044769f
C12342 a_11087_n20850.n49 VSS 0.129587f
C12343 a_11023_n4162.n0 VSS 0.016619f
C12344 a_11023_n4162.n1 VSS 0.646071f
C12345 a_11023_n4162.n2 VSS 0.0574f
C12346 a_11023_n4162.n3 VSS 0.016723f
C12347 a_11023_n4162.n4 VSS 0.057191f
C12348 a_11023_n4162.n5 VSS 0.056982f
C12349 a_11023_n4162.n6 VSS 0.056773f
C12350 a_11023_n4162.n7 VSS 0.318043f
C12351 a_11023_n4162.n8 VSS 0.318043f
C12352 a_11023_n4162.n9 VSS 0.318043f
C12353 a_11023_n4162.n10 VSS 0.440197f
C12354 a_11023_n4162.n11 VSS 0.107951f
C12355 a_11023_n4162.n12 VSS 0.052801f
C12356 a_11023_n4162.n13 VSS 0.022159f
C12357 a_11023_n4162.n14 VSS 0.052592f
C12358 a_11023_n4162.n15 VSS 0.022159f
C12359 a_11023_n4162.n16 VSS 0.052383f
C12360 a_11023_n4162.n17 VSS 0.052174f
C12361 a_11023_n4162.t15 VSS 0.038046f
C12362 a_11023_n4162.t17 VSS 0.038046f
C12363 a_11023_n4162.t11 VSS 0.038046f
C12364 a_11023_n4162.n18 VSS 0.198238f
C12365 a_11023_n4162.t37 VSS 0.064777f
C12366 a_11023_n4162.n19 VSS 0.145665f
C12367 a_11023_n4162.t30 VSS 0.06465f
C12368 a_11023_n4162.n20 VSS 0.056431f
C12369 a_11023_n4162.t34 VSS 0.06465f
C12370 a_11023_n4162.n21 VSS 0.016723f
C12371 a_11023_n4162.n22 VSS 0.120365f
C12372 a_11023_n4162.n23 VSS 0.022159f
C12373 a_11023_n4162.n24 VSS 0.022159f
C12374 a_11023_n4162.t39 VSS 0.06465f
C12375 a_11023_n4162.t28 VSS 0.06465f
C12376 a_11023_n4162.t23 VSS 0.06465f
C12377 a_11023_n4162.t35 VSS 0.06465f
C12378 a_11023_n4162.t36 VSS 0.064506f
C12379 a_11023_n4162.t25 VSS 0.064403f
C12380 a_11023_n4162.t21 VSS 0.064403f
C12381 a_11023_n4162.t38 VSS 0.064403f
C12382 a_11023_n4162.t27 VSS 0.064403f
C12383 a_11023_n4162.t22 VSS 0.064403f
C12384 a_11023_n4162.t32 VSS 0.064403f
C12385 a_11023_n4162.t24 VSS 0.064403f
C12386 a_11023_n4162.t20 VSS 0.064403f
C12387 a_11023_n4162.t29 VSS 0.064403f
C12388 a_11023_n4162.n25 VSS 0.223528f
C12389 a_11023_n4162.t26 VSS 0.06465f
C12390 a_11023_n4162.n26 VSS 0.072599f
C12391 a_11023_n4162.n27 VSS 0.022159f
C12392 a_11023_n4162.n28 VSS 0.016723f
C12393 a_11023_n4162.t31 VSS 0.06465f
C12394 a_11023_n4162.n29 VSS 0.022159f
C12395 a_11023_n4162.n30 VSS 0.022159f
C12396 a_11023_n4162.n31 VSS 0.016723f
C12397 a_11023_n4162.t33 VSS 0.06465f
C12398 a_11023_n4162.t6 VSS 0.038046f
C12399 a_11023_n4162.t4 VSS 0.038046f
C12400 a_11023_n4162.n32 VSS 0.180651f
C12401 a_11023_n4162.t3 VSS 0.038046f
C12402 a_11023_n4162.t0 VSS 0.038046f
C12403 a_11023_n4162.n33 VSS 0.180651f
C12404 a_11023_n4162.t2 VSS 0.038046f
C12405 a_11023_n4162.t8 VSS 0.038046f
C12406 a_11023_n4162.n34 VSS 0.180651f
C12407 a_11023_n4162.t9 VSS 0.038046f
C12408 a_11023_n4162.t5 VSS 0.038046f
C12409 a_11023_n4162.n35 VSS 0.180651f
C12410 a_11023_n4162.t7 VSS 0.038046f
C12411 a_11023_n4162.t1 VSS 0.038046f
C12412 a_11023_n4162.n36 VSS 0.200645f
C12413 a_11023_n4162.n37 VSS 0.702578f
C12414 a_11023_n4162.n38 VSS 0.300774f
C12415 a_11023_n4162.n39 VSS 0.300774f
C12416 a_11023_n4162.n40 VSS 0.418266f
C12417 a_11023_n4162.n41 VSS 0.725258f
C12418 a_11023_n4162.t16 VSS 0.038046f
C12419 a_11023_n4162.t14 VSS 0.038046f
C12420 a_11023_n4162.n42 VSS 0.183088f
C12421 a_11023_n4162.n43 VSS 0.322395f
C12422 a_11023_n4162.t13 VSS 0.038046f
C12423 a_11023_n4162.t10 VSS 0.038046f
C12424 a_11023_n4162.n44 VSS 0.183088f
C12425 a_11023_n4162.n45 VSS 0.186332f
C12426 a_11023_n4162.t12 VSS 0.038046f
C12427 a_11023_n4162.t18 VSS 0.038046f
C12428 a_11023_n4162.n46 VSS 0.183088f
C12429 a_11023_n4162.n47 VSS 0.186332f
C12430 a_11023_n4162.n48 VSS 0.507914f
C12431 a_11023_n4162.n49 VSS 0.183091f
C12432 a_11023_n4162.t19 VSS 0.038046f
C12433 a_29900_760.t1 VSS 0.12481f
C12434 a_29900_760.t0 VSS 0.076429f
C12435 a_29900_760.n0 VSS 0.304264f
C12436 a_29900_760.n1 VSS 0.304264f
C12437 a_29900_760.n2 VSS 0.638362f
C12438 a_29900_760.n3 VSS 0.919557f
C12439 a_29900_760.n4 VSS 1.46374f
C12440 a_29900_760.t14 VSS 0.080019f
C12441 a_29900_760.t17 VSS 0.070832f
C12442 a_29900_760.t12 VSS 0.081553f
C12443 a_29900_760.n5 VSS 0.096486f
C12444 a_29900_760.t3 VSS 0.087373f
C12445 a_29900_760.t8 VSS 0.081565f
C12446 a_29900_760.t13 VSS 0.087373f
C12447 a_29900_760.t10 VSS 0.070832f
C12448 a_29900_760.t16 VSS 0.081553f
C12449 a_29900_760.n6 VSS 0.093589f
C12450 a_29900_760.n7 VSS 1.36528f
C12451 a_29900_760.t15 VSS 0.079543f
C12452 a_29900_760.t6 VSS 0.081553f
C12453 a_29900_760.t2 VSS 0.070832f
C12454 a_29900_760.n8 VSS 0.096486f
C12455 a_29900_760.t7 VSS 0.087373f
C12456 a_29900_760.t11 VSS 0.081565f
C12457 a_29900_760.t5 VSS 0.087373f
C12458 a_29900_760.t4 VSS 0.070832f
C12459 a_29900_760.t9 VSS 0.081553f
C12460 a_29900_760.n9 VSS 0.093589f
C12461 a_29900_760.n10 VSS 0.241427f
C12462 a_29444_n4328.t3 VSS 0.153626f
C12463 a_29444_n4328.t2 VSS 0.153626f
C12464 a_29444_n4328.t1 VSS 0.153626f
C12465 a_29444_n4328.t0 VSS 0.21199f
C12466 a_29444_n4328.n0 VSS 1.7219f
C12467 a_29444_n4328.t5 VSS 0.104481f
C12468 a_29444_n4328.t6 VSS 0.155004f
C12469 a_29444_n4328.t8 VSS 0.060311f
C12470 a_29444_n4328.n1 VSS 0.390618f
C12471 a_29444_n4328.t9 VSS 0.174659f
C12472 a_29444_n4328.t7 VSS 0.142124f
C12473 a_29444_n4328.n2 VSS 2.27868f
C12474 a_29444_n4328.n3 VSS 4.38267f
C12475 a_29444_n4328.t4 VSS 0.116685f
C12476 a_22672_n2214.t1 VSS 0.073793f
C12477 a_22672_n2214.t2 VSS 0.044876f
C12478 a_22672_n2214.t0 VSS 0.013708f
C12479 a_22672_n2214.t3 VSS 0.053758f
C12480 a_22672_n2214.t4 VSS 0.026561f
C12481 a_22672_n2214.n0 VSS 0.820735f
C12482 a_22672_n2214.n1 VSS 1.16657f
C12483 a_22140_n6694.t1 VSS 0.105639f
C12484 a_22140_n6694.t0 VSS 0.014069f
C12485 a_22140_n6694.t17 VSS 0.021464f
C12486 a_22140_n6694.t13 VSS 0.016024f
C12487 a_22140_n6694.n0 VSS 0.107241f
C12488 a_22140_n6694.t16 VSS 0.010538f
C12489 a_22140_n6694.n1 VSS 0.059382f
C12490 a_22140_n6694.t6 VSS 0.010043f
C12491 a_22140_n6694.n2 VSS 0.038603f
C12492 a_22140_n6694.t8 VSS 0.024162f
C12493 a_22140_n6694.t4 VSS 0.014335f
C12494 a_22140_n6694.n3 VSS 0.030124f
C12495 a_22140_n6694.n4 VSS 0.151789f
C12496 a_22140_n6694.t3 VSS 0.024162f
C12497 a_22140_n6694.t15 VSS 0.014335f
C12498 a_22140_n6694.n5 VSS 0.043734f
C12499 a_22140_n6694.n6 VSS 0.204859f
C12500 a_22140_n6694.n7 VSS 0.321428f
C12501 a_22140_n6694.t5 VSS 0.018156f
C12502 a_22140_n6694.t2 VSS 0.023341f
C12503 a_22140_n6694.n8 VSS 0.036967f
C12504 a_22140_n6694.t9 VSS 0.010741f
C12505 a_22140_n6694.n9 VSS 0.052522f
C12506 a_22140_n6694.n10 VSS 0.299966f
C12507 a_22140_n6694.n11 VSS 0.420987f
C12508 a_22140_n6694.t10 VSS 0.010538f
C12509 a_22140_n6694.n12 VSS 0.03948f
C12510 a_22140_n6694.n13 VSS 0.332336f
C12511 a_22140_n6694.n14 VSS 0.404309f
C12512 a_25940_n17606.t1 VSS 0.085221f
C12513 a_25940_n17606.t0 VSS 0.044387f
C12514 a_25940_n17606.n0 VSS 0.934229f
C12515 a_25940_n17606.n1 VSS 0.503605f
C12516 a_25940_n17606.n2 VSS 1.2558f
C12517 a_25940_n17606.t7 VSS 0.045184f
C12518 a_25940_n17606.t9 VSS 0.047303f
C12519 a_25940_n17606.n3 VSS 0.055169f
C12520 a_25940_n17606.t23 VSS 0.022111f
C12521 a_25940_n17606.t14 VSS 0.020945f
C12522 a_25940_n17606.n4 VSS 0.154347f
C12523 a_25940_n17606.t4 VSS 0.020725f
C12524 a_25940_n17606.t25 VSS 0.022679f
C12525 a_25940_n17606.n5 VSS 0.062302f
C12526 a_25940_n17606.t11 VSS 0.041591f
C12527 a_25940_n17606.t6 VSS 0.048087f
C12528 a_25940_n17606.n6 VSS 0.078082f
C12529 a_25940_n17606.t22 VSS 0.041591f
C12530 a_25940_n17606.t2 VSS 0.048087f
C12531 a_25940_n17606.n7 VSS 0.07959f
C12532 a_25940_n17606.n8 VSS 0.699632f
C12533 a_25940_n17606.t18 VSS 0.023116f
C12534 a_25940_n17606.t17 VSS 0.020719f
C12535 a_25940_n17606.n9 VSS 0.058022f
C12536 a_25940_n17606.n10 VSS 0.661227f
C12537 a_25940_n17606.t15 VSS 0.041591f
C12538 a_25940_n17606.t3 VSS 0.048087f
C12539 a_25940_n17606.n11 VSS 0.079117f
C12540 a_25940_n17606.t10 VSS 0.023116f
C12541 a_25940_n17606.t12 VSS 0.020719f
C12542 a_25940_n17606.n12 VSS 0.060323f
C12543 a_25940_n17606.n13 VSS 0.206168f
C12544 a_25940_n17606.t20 VSS 0.023116f
C12545 a_25940_n17606.t21 VSS 0.020719f
C12546 a_25940_n17606.n14 VSS 0.057678f
C12547 a_25940_n17606.n15 VSS 0.174548f
C12548 a_25940_n17606.t19 VSS 0.041591f
C12549 a_25940_n17606.t8 VSS 0.048087f
C12550 a_25940_n17606.n16 VSS 0.111585f
C12551 a_25940_n17606.n17 VSS 0.981431f
C12552 a_25940_n17606.t5 VSS 0.04402f
C12553 a_25940_n17606.t13 VSS 0.044806f
C12554 a_25940_n17606.n18 VSS 0.069492f
C12555 a_25940_n17606.t24 VSS 0.023116f
C12556 a_25940_n17606.t16 VSS 0.020719f
C12557 a_25940_n17606.n19 VSS 0.058924f
C12558 a_25940_n17606.n20 VSS 0.42729f
C12559 a_32108_n2332.n0 VSS 0.437082f
C12560 a_32108_n2332.n1 VSS 0.18725f
C12561 a_32108_n2332.n2 VSS 0.130632f
C12562 a_32108_n2332.t14 VSS 0.027191f
C12563 a_32108_n2332.t13 VSS 0.027191f
C12564 a_32108_n2332.t11 VSS 0.027191f
C12565 a_32108_n2332.n3 VSS 0.067958f
C12566 a_32108_n2332.t9 VSS 0.027191f
C12567 a_32108_n2332.t12 VSS 0.027191f
C12568 a_32108_n2332.n4 VSS 0.055064f
C12569 a_32108_n2332.t10 VSS 0.027191f
C12570 a_32108_n2332.t8 VSS 0.027191f
C12571 a_32108_n2332.n5 VSS 0.055969f
C12572 a_32108_n2332.t21 VSS 0.035367f
C12573 a_32108_n2332.t23 VSS 0.039004f
C12574 a_32108_n2332.n6 VSS 0.090843f
C12575 a_32108_n2332.t17 VSS 0.039159f
C12576 a_32108_n2332.t18 VSS 0.035204f
C12577 a_32108_n2332.n7 VSS 0.081074f
C12578 a_32108_n2332.n8 VSS 0.44584f
C12579 a_32108_n2332.t16 VSS 0.039159f
C12580 a_32108_n2332.t20 VSS 0.035204f
C12581 a_32108_n2332.n9 VSS 0.096961f
C12582 a_32108_n2332.n10 VSS 0.843797f
C12583 a_32108_n2332.t22 VSS 0.039159f
C12584 a_32108_n2332.t24 VSS 0.035204f
C12585 a_32108_n2332.n11 VSS 0.078795f
C12586 a_32108_n2332.n12 VSS 0.526263f
C12587 a_32108_n2332.t26 VSS 0.035367f
C12588 a_32108_n2332.t27 VSS 0.039004f
C12589 a_32108_n2332.n13 VSS 0.255269f
C12590 a_32108_n2332.n14 VSS 0.790189f
C12591 a_32108_n2332.t25 VSS 0.035367f
C12592 a_32108_n2332.t19 VSS 0.039004f
C12593 a_32108_n2332.n15 VSS 0.081065f
C12594 a_32108_n2332.n16 VSS 0.434003f
C12595 a_32108_n2332.n17 VSS 0.014058f
C12596 a_32108_n2332.n18 VSS 0.019831f
C12597 a_32108_n2332.n19 VSS 0.014058f
C12598 a_32108_n2332.n20 VSS 0.019831f
C12599 a_32108_n2332.n21 VSS 0.055064f
C12600 a_32108_n2332.t15 VSS 0.027191f
C12601 a_35456_n4628.n0 VSS 0.466769f
C12602 a_35456_n4628.t4 VSS 0.024116f
C12603 a_35456_n4628.t0 VSS 0.021375f
C12604 a_35456_n4628.n1 VSS 0.025404f
C12605 a_35456_n4628.t13 VSS 0.076349f
C12606 a_35456_n4628.t17 VSS 0.04632f
C12607 a_35456_n4628.n2 VSS 0.111235f
C12608 a_35456_n4628.t18 VSS 0.076349f
C12609 a_35456_n4628.t15 VSS 0.04632f
C12610 a_35456_n4628.n3 VSS -0.029833f
C12611 a_35456_n4628.t11 VSS 0.076349f
C12612 a_35456_n4628.t16 VSS 0.04632f
C12613 a_35456_n4628.n4 VSS 0.126528f
C12614 a_35456_n4628.t12 VSS 0.076349f
C12615 a_35456_n4628.t9 VSS 0.04632f
C12616 a_35456_n4628.n5 VSS 0.126528f
C12617 a_35456_n4628.t20 VSS 0.076349f
C12618 a_35456_n4628.t8 VSS 0.04632f
C12619 a_35456_n4628.n6 VSS 0.126528f
C12620 a_35456_n4628.t14 VSS 0.076349f
C12621 a_35456_n4628.t10 VSS 0.04632f
C12622 a_35456_n4628.n7 VSS 0.12344f
C12623 a_35456_n4628.t22 VSS 0.076349f
C12624 a_35456_n4628.t21 VSS 0.04632f
C12625 a_35456_n4628.n8 VSS 0.111235f
C12626 a_35456_n4628.t19 VSS 0.076349f
C12627 a_35456_n4628.t7 VSS 0.04632f
C12628 a_35456_n4628.n9 VSS 0.114323f
C12629 a_35456_n4628.n10 VSS 0.074228f
C12630 a_35456_n4628.t5 VSS 0.024116f
C12631 a_35456_n4628.t3 VSS 0.024116f
C12632 a_35456_n4628.n11 VSS 0.058485f
C12633 a_35456_n4628.n12 VSS 0.04873f
C12634 a_35456_n4628.t6 VSS 0.024116f
C12635 a_28736_n4633.n0 VSS 0.453203f
C12636 a_28736_n4633.n1 VSS 0.392182f
C12637 a_28736_n4633.n2 VSS 0.398956f
C12638 a_28736_n4633.t10 VSS 0.018674f
C12639 a_28736_n4633.t16 VSS 0.033456f
C12640 a_28736_n4633.t15 VSS 0.033456f
C12641 a_28736_n4633.n3 VSS 0.080174f
C12642 a_28736_n4633.t14 VSS 0.033456f
C12643 a_28736_n4633.t17 VSS 0.033456f
C12644 a_28736_n4633.n4 VSS 0.059261f
C12645 a_28736_n4633.n5 VSS 0.25634f
C12646 a_28736_n4633.t12 VSS 0.018674f
C12647 a_28736_n4633.t0 VSS 0.018674f
C12648 a_28736_n4633.n6 VSS 0.037885f
C12649 a_28736_n4633.t1 VSS 0.018674f
C12650 a_28736_n4633.t13 VSS 0.018674f
C12651 a_28736_n4633.n7 VSS 0.037885f
C12652 a_28736_n4633.t11 VSS 0.018674f
C12653 a_28736_n4633.t2 VSS 0.018674f
C12654 a_28736_n4633.n8 VSS 0.037885f
C12655 a_28736_n4633.t8 VSS 0.018674f
C12656 a_28736_n4633.t5 VSS 0.018674f
C12657 a_28736_n4633.n9 VSS 0.037885f
C12658 a_28736_n4633.t4 VSS 0.018674f
C12659 a_28736_n4633.t9 VSS 0.018674f
C12660 a_28736_n4633.n10 VSS 0.037885f
C12661 a_28736_n4633.t7 VSS 0.018674f
C12662 a_28736_n4633.t6 VSS 0.018674f
C12663 a_28736_n4633.n11 VSS 0.037885f
C12664 a_28736_n4633.t19 VSS 0.018674f
C12665 a_28736_n4633.t18 VSS 0.018674f
C12666 a_28736_n4633.n12 VSS 0.04653f
C12667 a_28736_n4633.t21 VSS 0.084749f
C12668 a_28736_n4633.t25 VSS 0.085142f
C12669 a_28736_n4633.t20 VSS 0.073949f
C12670 a_28736_n4633.n13 VSS 0.100732f
C12671 a_28736_n4633.t22 VSS 0.091218f
C12672 a_28736_n4633.t24 VSS 0.070025f
C12673 a_28736_n4633.t23 VSS 0.080961f
C12674 a_28736_n4633.n14 VSS 0.736029f
C12675 a_28736_n4633.n15 VSS 1.59544f
C12676 a_28736_n4633.n16 VSS 0.197307f
C12677 a_28736_n4633.n17 VSS 0.037885f
C12678 a_28736_n4633.t3 VSS 0.018674f
C12679 a_30452_n5156.n0 VSS 0.504151f
C12680 a_30452_n5156.t2 VSS 0.110214f
C12681 a_30452_n5156.n1 VSS 0.024426f
C12682 a_30452_n5156.t9 VSS 0.067227f
C12683 a_30452_n5156.t5 VSS 0.063923f
C12684 a_30452_n5156.n2 VSS 0.099029f
C12685 a_30452_n5156.t10 VSS 0.067227f
C12686 a_30452_n5156.t4 VSS 0.063923f
C12687 a_30452_n5156.n3 VSS 0.096963f
C12688 a_30452_n5156.n4 VSS 0.071087f
C12689 a_30452_n5156.t7 VSS 0.052924f
C12690 a_30452_n5156.n5 VSS 0.044088f
C12691 a_30452_n5156.t14 VSS 0.06134f
C12692 a_30452_n5156.n6 VSS 0.072876f
C12693 a_30452_n5156.t6 VSS 0.06134f
C12694 a_30452_n5156.n7 VSS 0.072876f
C12695 a_30452_n5156.t11 VSS 0.052924f
C12696 a_30452_n5156.n8 VSS 0.042206f
C12697 a_30452_n5156.t8 VSS 0.06134f
C12698 a_30452_n5156.t3 VSS 0.06134f
C12699 a_30452_n5156.t12 VSS 0.052924f
C12700 a_30452_n5156.n9 VSS 0.042206f
C12701 a_30452_n5156.n10 VSS 0.072876f
C12702 a_30452_n5156.n11 VSS 0.072876f
C12703 a_30452_n5156.t13 VSS 0.052924f
C12704 a_30452_n5156.n12 VSS 0.042206f
C12705 a_30452_n5156.n13 VSS 1.26513f
C12706 a_30452_n5156.n14 VSS 0.729337f
C12707 a_21692_n13308.n0 VSS 0.349631f
C12708 a_21692_n13308.n1 VSS 0.522674f
C12709 a_21692_n13308.n2 VSS 0.290887f
C12710 a_21692_n13308.t10 VSS 0.029907f
C12711 a_21692_n13308.t14 VSS 0.029907f
C12712 a_21692_n13308.t13 VSS 0.029907f
C12713 a_21692_n13308.n3 VSS 0.074746f
C12714 a_21692_n13308.t11 VSS 0.029907f
C12715 a_21692_n13308.t8 VSS 0.029907f
C12716 a_21692_n13308.n4 VSS 0.060563f
C12717 a_21692_n13308.t12 VSS 0.029907f
C12718 a_21692_n13308.t9 VSS 0.029907f
C12719 a_21692_n13308.n5 VSS 0.067638f
C12720 a_21692_n13308.t17 VSS 0.0389f
C12721 a_21692_n13308.t26 VSS 0.042899f
C12722 a_21692_n13308.n6 VSS 0.086655f
C12723 a_21692_n13308.t20 VSS 0.04307f
C12724 a_21692_n13308.t21 VSS 0.03872f
C12725 a_21692_n13308.n7 VSS 0.138994f
C12726 a_21692_n13308.t23 VSS 0.04307f
C12727 a_21692_n13308.t18 VSS 0.03872f
C12728 a_21692_n13308.n8 VSS 0.086482f
C12729 a_21692_n13308.n9 VSS 0.878451f
C12730 a_21692_n13308.t25 VSS 0.04307f
C12731 a_21692_n13308.t22 VSS 0.03872f
C12732 a_21692_n13308.n10 VSS 0.106645f
C12733 a_21692_n13308.n11 VSS 0.933653f
C12734 a_21692_n13308.t30 VSS 0.0389f
C12735 a_21692_n13308.t24 VSS 0.042899f
C12736 a_21692_n13308.n12 VSS 0.145754f
C12737 a_21692_n13308.n13 VSS 0.690299f
C12738 a_21692_n13308.t27 VSS 0.0389f
C12739 a_21692_n13308.t31 VSS 0.042899f
C12740 a_21692_n13308.n14 VSS 0.087425f
C12741 a_21692_n13308.n15 VSS 0.385068f
C12742 a_21692_n13308.t29 VSS 0.0389f
C12743 a_21692_n13308.t16 VSS 0.042899f
C12744 a_21692_n13308.n16 VSS 0.089162f
C12745 a_21692_n13308.n17 VSS 0.356789f
C12746 a_21692_n13308.t28 VSS 0.0389f
C12747 a_21692_n13308.t32 VSS 0.042899f
C12748 a_21692_n13308.n18 VSS 0.086655f
C12749 a_21692_n13308.n19 VSS 0.34986f
C12750 a_21692_n13308.t19 VSS 0.0389f
C12751 a_21692_n13308.t33 VSS 0.042899f
C12752 a_21692_n13308.n20 VSS 0.086655f
C12753 a_21692_n13308.n21 VSS 0.38269f
C12754 a_21692_n13308.n22 VSS 0.87119f
C12755 a_21692_n13308.n23 VSS 0.015463f
C12756 a_21692_n13308.n24 VSS 0.021812f
C12757 a_21692_n13308.n25 VSS 0.015463f
C12758 a_21692_n13308.n26 VSS 0.021812f
C12759 a_21692_n13308.n27 VSS 0.060563f
C12760 a_21692_n13308.t15 VSS 0.029907f
C12761 a_26328_n6654.n0 VSS 0.466769f
C12762 a_26328_n6654.t5 VSS 0.024116f
C12763 a_26328_n6654.t4 VSS 0.024116f
C12764 a_26328_n6654.t3 VSS 0.024116f
C12765 a_26328_n6654.n1 VSS 0.058485f
C12766 a_26328_n6654.t1 VSS 0.021375f
C12767 a_26328_n6654.n2 VSS 0.025404f
C12768 a_26328_n6654.t10 VSS 0.076349f
C12769 a_26328_n6654.t18 VSS 0.04632f
C12770 a_26328_n6654.n3 VSS 0.111235f
C12771 a_26328_n6654.t11 VSS 0.076349f
C12772 a_26328_n6654.t15 VSS 0.04632f
C12773 a_26328_n6654.n4 VSS 0.114323f
C12774 a_26328_n6654.t20 VSS 0.076349f
C12775 a_26328_n6654.t7 VSS 0.04632f
C12776 a_26328_n6654.n5 VSS 0.111235f
C12777 a_26328_n6654.t13 VSS 0.076349f
C12778 a_26328_n6654.t22 VSS 0.04632f
C12779 a_26328_n6654.n6 VSS -0.029833f
C12780 a_26328_n6654.t21 VSS 0.076349f
C12781 a_26328_n6654.t8 VSS 0.04632f
C12782 a_26328_n6654.n7 VSS 0.126528f
C12783 a_26328_n6654.t16 VSS 0.076349f
C12784 a_26328_n6654.t12 VSS 0.04632f
C12785 a_26328_n6654.n8 VSS 0.126528f
C12786 a_26328_n6654.t9 VSS 0.076349f
C12787 a_26328_n6654.t14 VSS 0.04632f
C12788 a_26328_n6654.n9 VSS 0.126528f
C12789 a_26328_n6654.t19 VSS 0.076349f
C12790 a_26328_n6654.t17 VSS 0.04632f
C12791 a_26328_n6654.n10 VSS 0.12344f
C12792 a_26328_n6654.n11 VSS 0.074228f
C12793 a_26328_n6654.n12 VSS 0.04873f
C12794 a_26328_n6654.t6 VSS 0.024116f
C12795 a_24481_761.n0 VSS 0.395705f
C12796 a_24481_761.n1 VSS 0.297312f
C12797 a_24481_761.n2 VSS 0.350459f
C12798 a_24481_761.t6 VSS 0.025297f
C12799 a_24481_761.t5 VSS 0.020961f
C12800 a_24481_761.t4 VSS 0.020961f
C12801 a_24481_761.t7 VSS 0.025297f
C12802 a_24481_761.n3 VSS 0.600186f
C12803 a_24481_761.n4 VSS 0.499558f
C12804 a_24481_761.n5 VSS 0.500916f
C12805 a_24481_761.n6 VSS 0.426699f
C12806 a_24481_761.n7 VSS 0.439748f
C12807 a_24481_761.t0 VSS 0.091906f
C12808 a_24481_761.n8 VSS 0.597487f
C12809 a_24481_761.n9 VSS 0.057964f
C12810 a_24481_761.n10 VSS 0.825854f
C12811 a_24481_761.t1 VSS 0.056256f
C12812 a_24481_761.n11 VSS 0.41959f
C12813 a_24481_761.t3 VSS 0.055522f
C12814 a_24481_761.t2 VSS 0.055522f
C12815 a_24481_761.t42 VSS 0.019093f
C12816 a_24481_761.t47 VSS 0.020892f
C12817 a_24481_761.n12 VSS 0.066162f
C12818 a_24481_761.t59 VSS 0.021295f
C12819 a_24481_761.t85 VSS 0.019087f
C12820 a_24481_761.n13 VSS 0.067488f
C12821 a_24481_761.t19 VSS 0.019296f
C12822 a_24481_761.t10 VSS 0.02037f
C12823 a_24481_761.n14 VSS 0.084541f
C12824 a_24481_761.t44 VSS 0.021295f
C12825 a_24481_761.t63 VSS 0.019087f
C12826 a_24481_761.n15 VSS 0.07792f
C12827 a_24481_761.t84 VSS 0.057902f
C12828 a_24481_761.t14 VSS 0.055286f
C12829 a_24481_761.t87 VSS 0.162609f
C12830 a_24481_761.t93 VSS 0.122156f
C12831 a_24481_761.n16 VSS 0.079485f
C12832 a_24481_761.t56 VSS 0.057902f
C12833 a_24481_761.t67 VSS 0.055286f
C12834 a_24481_761.t22 VSS 0.162609f
C12835 a_24481_761.t8 VSS 0.122156f
C12836 a_24481_761.n17 VSS 0.103067f
C12837 a_24481_761.t78 VSS 0.027289f
C12838 a_24481_761.t50 VSS 0.060153f
C12839 a_24481_761.t45 VSS 0.139014f
C12840 a_24481_761.t82 VSS 0.107644f
C12841 a_24481_761.n18 VSS 0.060378f
C12842 a_24481_761.n19 VSS 0.500336f
C12843 a_24481_761.t58 VSS 0.057902f
C12844 a_24481_761.t27 VSS 0.055286f
C12845 a_24481_761.t89 VSS 0.162609f
C12846 a_24481_761.t80 VSS 0.120706f
C12847 a_24481_761.n20 VSS 0.089861f
C12848 a_24481_761.t17 VSS 0.020892f
C12849 a_24481_761.t48 VSS 0.019093f
C12850 a_24481_761.t92 VSS 0.020892f
C12851 a_24481_761.t36 VSS 0.019093f
C12852 a_24481_761.n21 VSS 0.061562f
C12853 a_24481_761.n22 VSS 0.690761f
C12854 a_24481_761.t57 VSS 0.021295f
C12855 a_24481_761.t83 VSS 0.019087f
C12856 a_24481_761.n23 VSS 0.054284f
C12857 a_24481_761.t86 VSS 0.057902f
C12858 a_24481_761.t66 VSS 0.055286f
C12859 a_24481_761.t31 VSS 0.162609f
C12860 a_24481_761.t46 VSS 0.122156f
C12861 a_24481_761.n24 VSS 0.059334f
C12862 a_24481_761.t24 VSS 0.021295f
C12863 a_24481_761.t43 VSS 0.019087f
C12864 a_24481_761.n25 VSS 0.053135f
C12865 a_24481_761.t16 VSS 0.021295f
C12866 a_24481_761.t52 VSS 0.019087f
C12867 a_24481_761.n26 VSS 0.053436f
C12868 a_24481_761.t21 VSS 0.055286f
C12869 a_24481_761.t61 VSS 0.162609f
C12870 a_24481_761.t12 VSS 0.122156f
C12871 a_24481_761.t54 VSS 0.057902f
C12872 a_24481_761.n27 VSS 0.083408f
C12873 a_24481_761.t49 VSS 0.057902f
C12874 a_24481_761.t81 VSS 0.055286f
C12875 a_24481_761.t51 VSS 0.162609f
C12876 a_24481_761.t71 VSS 0.122156f
C12877 a_24481_761.n28 VSS 0.159952f
C12878 a_24481_761.t53 VSS 0.021295f
C12879 a_24481_761.t79 VSS 0.019087f
C12880 a_24481_761.n29 VSS 0.053135f
C12881 a_24481_761.n30 VSS 0.35742f
C12882 a_24481_761.t65 VSS 0.021295f
C12883 a_24481_761.t55 VSS 0.019087f
C12884 a_24481_761.n31 VSS 0.135977f
C12885 a_24481_761.n32 VSS 0.460972f
C12886 a_24481_761.t11 VSS 0.057902f
C12887 a_24481_761.t60 VSS 0.055286f
C12888 a_24481_761.t28 VSS 0.162609f
C12889 a_24481_761.t70 VSS 0.122156f
C12890 a_24481_761.n33 VSS 0.052021f
C12891 a_24481_761.t90 VSS 0.055286f
C12892 a_24481_761.t35 VSS 0.162609f
C12893 a_24481_761.t68 VSS 0.122156f
C12894 a_24481_761.t18 VSS 0.059715f
C12895 a_24481_761.n34 VSS 0.184833f
C12896 a_24481_761.t34 VSS 0.021295f
C12897 a_24481_761.t76 VSS 0.019087f
C12898 a_24481_761.n35 VSS 0.053135f
C12899 a_24481_761.t72 VSS 0.057902f
C12900 a_24481_761.t62 VSS 0.055286f
C12901 a_24481_761.t29 VSS 0.162609f
C12902 a_24481_761.t33 VSS 0.122156f
C12903 a_24481_761.n36 VSS 0.051904f
C12904 a_24481_761.n37 VSS 0.235337f
C12905 a_24481_761.t9 VSS 0.055286f
C12906 a_24481_761.t94 VSS 0.162609f
C12907 a_24481_761.t15 VSS 0.122156f
C12908 a_24481_761.t13 VSS 0.059715f
C12909 a_24481_761.n38 VSS 0.102694f
C12910 a_24481_761.t64 VSS 0.055286f
C12911 a_24481_761.t77 VSS 0.162609f
C12912 a_24481_761.t73 VSS 0.122156f
C12913 a_24481_761.t38 VSS 0.057902f
C12914 a_24481_761.n39 VSS 0.057896f
C12915 a_24481_761.n40 VSS 0.678877f
C12916 a_24481_761.t75 VSS 0.019912f
C12917 a_24481_761.t69 VSS 0.019504f
C12918 a_24481_761.n41 VSS 0.305f
C12919 a_24481_761.t32 VSS 0.055286f
C12920 a_24481_761.t30 VSS 0.162609f
C12921 a_24481_761.t39 VSS 0.122156f
C12922 a_24481_761.t41 VSS 0.057902f
C12923 a_24481_761.n42 VSS 0.117063f
C12924 a_24481_761.n43 VSS 0.657915f
C12925 a_24481_761.t74 VSS 0.05882f
C12926 a_24481_761.t23 VSS 0.038782f
C12927 a_24481_761.t37 VSS 0.021766f
C12928 a_24481_761.n44 VSS 0.103763f
C12929 a_24481_761.t26 VSS 0.038782f
C12930 a_24481_761.t40 VSS 0.021766f
C12931 a_24481_761.n45 VSS 0.067035f
C12932 a_24481_761.t88 VSS 0.038782f
C12933 a_24481_761.t20 VSS 0.021766f
C12934 a_24481_761.t25 VSS 0.019093f
C12935 a_24481_761.t91 VSS 0.020892f
C12936 a_24481_761.n46 VSS 0.602447f
C12937 a_13501_n22528.n0 VSS 2.0189f
C12938 a_13501_n22528.n1 VSS 3.79312f
C12939 a_13501_n22528.t15 VSS 0.041646f
C12940 a_13501_n22528.t11 VSS 0.33153f
C12941 a_13501_n22528.t2 VSS 0.321965f
C12942 a_13501_n22528.t0 VSS 0.041646f
C12943 a_13501_n22528.t4 VSS 0.041646f
C12944 a_13501_n22528.n2 VSS 0.229216f
C12945 a_13501_n22528.t19 VSS 0.041646f
C12946 a_13501_n22528.t13 VSS 0.041646f
C12947 a_13501_n22528.n3 VSS 0.223712f
C12948 a_13501_n22528.t7 VSS 0.041646f
C12949 a_13501_n22528.t1 VSS 0.041646f
C12950 a_13501_n22528.n4 VSS 0.228449f
C12951 a_13501_n22528.t16 VSS 0.041646f
C12952 a_13501_n22528.t10 VSS 0.041646f
C12953 a_13501_n22528.n5 VSS 0.22515f
C12954 a_13501_n22528.t14 VSS 0.041646f
C12955 a_13501_n22528.t17 VSS 0.041646f
C12956 a_13501_n22528.n6 VSS 0.22515f
C12957 a_13501_n22528.t5 VSS 0.041646f
C12958 a_13501_n22528.t8 VSS 0.041646f
C12959 a_13501_n22528.n7 VSS 0.227874f
C12960 a_13501_n22528.t6 VSS 0.041646f
C12961 a_13501_n22528.t9 VSS 0.041646f
C12962 a_13501_n22528.n8 VSS 0.228065f
C12963 a_13501_n22528.t12 VSS 0.33124f
C12964 a_13501_n22528.t3 VSS 0.325425f
C12965 a_13501_n22528.n9 VSS 0.22387f
C12966 a_13501_n22528.t18 VSS 0.041646f
C12967 a_21692_n5111.t0 VSS 0.010486f
C12968 a_21692_n5111.t3 VSS 0.031124f
C12969 a_21692_n5111.t2 VSS 0.016396f
C12970 a_21692_n5111.n0 VSS 0.24669f
C12971 a_21692_n5111.t4 VSS 0.031124f
C12972 a_21692_n5111.t5 VSS 0.016396f
C12973 a_21692_n5111.n1 VSS 0.033163f
C12974 a_21692_n5111.n2 VSS 1.15508f
C12975 a_21692_n5111.n3 VSS 0.430237f
C12976 a_21692_n5111.t1 VSS 0.029302f
C12977 OUT[3].t13 VSS 0.030992f
C12978 OUT[3].t11 VSS 0.022383f
C12979 OUT[3].n0 VSS 0.054045f
C12980 OUT[3].t8 VSS 0.030992f
C12981 OUT[3].t14 VSS 0.022383f
C12982 OUT[3].n1 VSS 0.054045f
C12983 OUT[3].t12 VSS 0.030992f
C12984 OUT[3].t10 VSS 0.022383f
C12985 OUT[3].n2 VSS 0.068367f
C12986 OUT[3].n3 VSS 0.172904f
C12987 OUT[3].t6 VSS 0.015044f
C12988 OUT[3].t4 VSS 0.015044f
C12989 OUT[3].n4 VSS 0.030193f
C12990 OUT[3].t2 VSS 0.015044f
C12991 OUT[3].t0 VSS 0.015044f
C12992 OUT[3].n5 VSS 0.036302f
C12993 OUT[3].n6 VSS 0.162383f
C12994 OUT[3].t1 VSS 0.015044f
C12995 OUT[3].t7 VSS 0.015044f
C12996 OUT[3].n7 VSS 0.030193f
C12997 OUT[3].t5 VSS 0.015044f
C12998 OUT[3].t3 VSS 0.015044f
C12999 OUT[3].n8 VSS 0.036182f
C13000 OUT[3].n9 VSS 0.165248f
C13001 OUT[3].n10 VSS 0.132888f
C13002 OUT[3].n11 VSS 0.132888f
C13003 OUT[3].n12 VSS 0.108893f
C13004 OUT[3].t9 VSS 0.022383f
C13005 OUT[3].t15 VSS 0.030992f
C13006 OUT[3].n13 VSS 0.053376f
C13007 OUT[3].n14 VSS 0.396132f
C13008 a_22220_690.n0 VSS 0.105728f
C13009 a_22220_690.n1 VSS 2.79321f
C13010 a_22220_690.t1 VSS 0.32041f
C13011 a_22220_690.n2 VSS 3.46796f
C13012 a_22220_690.t0 VSS 0.053452f
C13013 a_22220_690.t11 VSS 0.039228f
C13014 a_22220_690.t13 VSS 0.035161f
C13015 a_22220_690.n3 VSS 0.68398f
C13016 a_22220_690.t10 VSS 0.038486f
C13017 a_22220_690.t5 VSS 0.035172f
C13018 a_22220_690.t16 VSS 0.085247f
C13019 a_22220_690.t14 VSS 0.066308f
C13020 a_22220_690.n4 VSS 0.152544f
C13021 a_22220_690.t7 VSS 0.079767f
C13022 a_22220_690.t9 VSS 0.067469f
C13023 a_22220_690.n5 VSS 0.182243f
C13024 a_22220_690.t12 VSS 0.069654f
C13025 a_22220_690.t8 VSS 0.085599f
C13026 a_22220_690.n6 VSS 0.828639f
C13027 a_22220_690.t15 VSS 0.039228f
C13028 a_22220_690.t6 VSS 0.035161f
C13029 a_22220_690.n7 VSS 0.09788f
C13030 a_22220_690.n8 VSS 1.87342f
C13031 a_22220_690.t17 VSS 0.067832f
C13032 a_22220_690.t2 VSS 0.077964f
C13033 a_22220_690.n9 VSS 0.127408f
C13034 a_22220_690.n10 VSS 1.81276f
C13035 a_22220_690.t4 VSS 0.036681f
C13036 a_22220_690.t3 VSS 0.035929f
C13037 a_22220_690.n11 VSS 0.119251f
C13038 a_22220_690.n12 VSS 0.686232f
C13039 a_28519_n10160.t1 VSS 0.424247f
C13040 a_28519_n10160.t0 VSS 0.048928f
C13041 a_28519_n10160.t8 VSS 0.080768f
C13042 a_28519_n10160.t4 VSS 0.043926f
C13043 a_28519_n10160.n0 VSS 0.161203f
C13044 a_28519_n10160.t2 VSS 0.081991f
C13045 a_28519_n10160.t7 VSS 0.061677f
C13046 a_28519_n10160.n1 VSS 0.097907f
C13047 a_28519_n10160.t3 VSS 0.062811f
C13048 a_28519_n10160.t5 VSS 0.085255f
C13049 a_28519_n10160.n2 VSS 0.129454f
C13050 a_28519_n10160.n3 VSS 0.97982f
C13051 a_28519_n10160.t9 VSS 0.079648f
C13052 a_28519_n10160.t6 VSS 0.069754f
C13053 a_28519_n10160.n4 VSS 0.176068f
C13054 a_28519_n10160.n5 VSS 1.21654f
C13055 a_25612_n878.n0 VSS 0.111339f
C13056 a_25612_n878.t0 VSS 0.039991f
C13057 a_25612_n878.t1 VSS 0.022537f
C13058 a_25612_n878.t3 VSS 0.029084f
C13059 a_25612_n878.t4 VSS 0.037391f
C13060 a_25612_n878.n1 VSS 0.099702f
C13061 a_25612_n878.t5 VSS 0.030552f
C13062 a_25612_n878.t6 VSS 0.037546f
C13063 a_25612_n878.n2 VSS 0.118286f
C13064 a_25612_n878.t2 VSS 0.038707f
C13065 a_25612_n878.t7 VSS 0.022964f
C13066 a_25612_n878.n3 VSS 0.078323f
C13067 a_25612_n878.n4 VSS 0.895886f
C13068 a_25612_n878.n5 VSS 0.737691f
C13069 a_27259_804.n0 VSS 1.0865f
C13070 a_27259_804.n1 VSS 0.14825f
C13071 a_27259_804.t0 VSS 0.060015f
C13072 a_27259_804.t1 VSS 0.070481f
C13073 a_27259_804.n2 VSS 1.41575f
C13074 a_27259_804.t2 VSS 0.044499f
C13075 a_27259_804.t13 VSS 0.057208f
C13076 a_27259_804.n3 VSS 0.342285f
C13077 a_27259_804.t5 VSS 0.045521f
C13078 a_27259_804.t4 VSS 0.052321f
C13079 a_27259_804.n4 VSS 0.301693f
C13080 a_27259_804.t6 VSS 0.039438f
C13081 a_27259_804.t12 VSS 0.052609f
C13082 a_27259_804.n5 VSS 0.090338f
C13083 a_27259_804.t16 VSS 0.041052f
C13084 a_27259_804.t3 VSS 0.052095f
C13085 a_27259_804.t14 VSS 0.049015f
C13086 a_27259_804.n6 VSS 0.076874f
C13087 a_27259_804.t19 VSS 0.048554f
C13088 a_27259_804.t15 VSS 0.04755f
C13089 a_27259_804.t8 VSS 0.054851f
C13090 a_27259_804.n7 VSS 0.096626f
C13091 a_27259_804.t11 VSS 0.048153f
C13092 a_27259_804.t9 VSS 0.055428f
C13093 a_27259_804.n8 VSS 0.087397f
C13094 a_27259_804.t7 VSS 0.04755f
C13095 a_27259_804.t18 VSS 0.054851f
C13096 a_27259_804.n9 VSS 0.107389f
C13097 a_27259_804.t17 VSS 0.04755f
C13098 a_27259_804.t10 VSS 0.054851f
C13099 a_27259_804.n10 VSS 0.223302f
C13100 a_21772_n452.n0 VSS 0.588053f
C13101 a_21772_n452.t2 VSS 0.052911f
C13102 a_21772_n452.t3 VSS 0.058323f
C13103 a_21772_n452.t0 VSS 0.07776f
C13104 a_21772_n452.t1 VSS 0.065058f
C13105 a_21772_n452.t7 VSS 0.058056f
C13106 a_21772_n452.t18 VSS 0.055202f
C13107 a_21772_n452.n1 VSS 0.090091f
C13108 a_21772_n452.t8 VSS 0.058056f
C13109 a_21772_n452.t12 VSS 0.055202f
C13110 a_21772_n452.n2 VSS 0.090091f
C13111 a_21772_n452.t6 VSS 0.058056f
C13112 a_21772_n452.t10 VSS 0.055202f
C13113 a_21772_n452.n3 VSS -0.035108f
C13114 a_21772_n452.t9 VSS 0.058056f
C13115 a_21772_n452.t17 VSS 0.055202f
C13116 a_21772_n452.n4 VSS 0.101689f
C13117 a_21772_n452.t5 VSS 0.058056f
C13118 a_21772_n452.t13 VSS 0.055202f
C13119 a_21772_n452.n5 VSS 0.101689f
C13120 a_21772_n452.t15 VSS 0.058056f
C13121 a_21772_n452.t11 VSS 0.055202f
C13122 a_21772_n452.n6 VSS 0.101689f
C13123 a_21772_n452.t4 VSS 0.058056f
C13124 a_21772_n452.t16 VSS 0.055202f
C13125 a_21772_n452.n7 VSS 0.101689f
C13126 a_21772_n452.t19 VSS 0.058056f
C13127 a_21772_n452.t14 VSS 0.055202f
C13128 a_30732_332.t1 VSS 0.536403f
C13129 a_30732_332.t3 VSS 0.016959f
C13130 a_30732_332.t5 VSS 0.034324f
C13131 a_30732_332.n0 VSS 0.272513f
C13132 a_30732_332.t7 VSS 0.018458f
C13133 a_30732_332.t2 VSS 0.035039f
C13134 a_30732_332.n1 VSS 0.075764f
C13135 a_30732_332.n2 VSS 0.740998f
C13136 a_30732_332.t4 VSS 0.029605f
C13137 a_30732_332.t6 VSS 0.035313f
C13138 a_30732_332.n3 VSS 0.18098f
C13139 a_30732_332.t0 VSS 0.023644f
C13140 a_13501_n11816.n0 VSS 2.0189f
C13141 a_13501_n11816.n1 VSS 3.79312f
C13142 a_13501_n11816.t2 VSS 0.041646f
C13143 a_13501_n11816.t5 VSS 0.33153f
C13144 a_13501_n11816.t13 VSS 0.321965f
C13145 a_13501_n11816.t15 VSS 0.041646f
C13146 a_13501_n11816.t11 VSS 0.041646f
C13147 a_13501_n11816.n2 VSS 0.229216f
C13148 a_13501_n11816.t3 VSS 0.041646f
C13149 a_13501_n11816.t7 VSS 0.041646f
C13150 a_13501_n11816.n3 VSS 0.223712f
C13151 a_13501_n11816.t18 VSS 0.041646f
C13152 a_13501_n11816.t14 VSS 0.041646f
C13153 a_13501_n11816.n4 VSS 0.228449f
C13154 a_13501_n11816.t0 VSS 0.041646f
C13155 a_13501_n11816.t4 VSS 0.041646f
C13156 a_13501_n11816.n5 VSS 0.22515f
C13157 a_13501_n11816.t8 VSS 0.041646f
C13158 a_13501_n11816.t1 VSS 0.041646f
C13159 a_13501_n11816.n6 VSS 0.22515f
C13160 a_13501_n11816.t10 VSS 0.041646f
C13161 a_13501_n11816.t17 VSS 0.041646f
C13162 a_13501_n11816.n7 VSS 0.227874f
C13163 a_13501_n11816.t19 VSS 0.041646f
C13164 a_13501_n11816.t16 VSS 0.041646f
C13165 a_13501_n11816.n8 VSS 0.228065f
C13166 a_13501_n11816.t6 VSS 0.33124f
C13167 a_13501_n11816.t12 VSS 0.325425f
C13168 a_13501_n11816.n9 VSS 0.22387f
C13169 a_13501_n11816.t9 VSS 0.041646f
C13170 a_31548_n10172.n0 VSS 0.468001f
C13171 a_31548_n10172.n1 VSS 0.082474f
C13172 a_31548_n10172.n2 VSS 0.132096f
C13173 a_31548_n10172.t10 VSS 0.027496f
C13174 a_31548_n10172.t12 VSS 0.027496f
C13175 a_31548_n10172.t11 VSS 0.027496f
C13176 a_31548_n10172.n3 VSS 0.05568f
C13177 a_31548_n10172.t13 VSS 0.027496f
C13178 a_31548_n10172.t9 VSS 0.027496f
C13179 a_31548_n10172.n4 VSS 0.068719f
C13180 a_31548_n10172.n5 VSS 0.014216f
C13181 a_31548_n10172.n6 VSS 0.020053f
C13182 a_31548_n10172.n7 VSS 0.014216f
C13183 a_31548_n10172.n8 VSS 0.020053f
C13184 a_31548_n10172.t8 VSS 0.027496f
C13185 a_31548_n10172.t14 VSS 0.027496f
C13186 a_31548_n10172.n9 VSS 0.058874f
C13187 a_31548_n10172.t22 VSS 0.039597f
C13188 a_31548_n10172.t19 VSS 0.035598f
C13189 a_31548_n10172.n10 VSS 0.171188f
C13190 a_31548_n10172.t17 VSS 0.039597f
C13191 a_31548_n10172.t24 VSS 0.035598f
C13192 a_31548_n10172.n11 VSS 0.153288f
C13193 a_31548_n10172.n12 VSS 0.742789f
C13194 a_31548_n10172.t16 VSS 0.035764f
C13195 a_31548_n10172.t25 VSS 0.039441f
C13196 a_31548_n10172.n13 VSS 0.155857f
C13197 a_31548_n10172.n14 VSS 0.311042f
C13198 a_31548_n10172.t18 VSS 0.035764f
C13199 a_31548_n10172.t23 VSS 0.039441f
C13200 a_31548_n10172.n15 VSS 0.174442f
C13201 a_31548_n10172.t20 VSS 0.035764f
C13202 a_31548_n10172.t21 VSS 0.039441f
C13203 a_31548_n10172.n16 VSS 0.221514f
C13204 a_31548_n10172.n17 VSS 1.11255f
C13205 a_31548_n10172.n18 VSS 0.315306f
C13206 a_31548_n10172.n19 VSS 0.05568f
C13207 a_31548_n10172.t15 VSS 0.027496f
C13208 a_33496_n8222.n0 VSS 0.466769f
C13209 a_33496_n8222.t4 VSS 0.024116f
C13210 a_33496_n8222.t3 VSS 0.024116f
C13211 a_33496_n8222.t5 VSS 0.024116f
C13212 a_33496_n8222.n1 VSS 0.04873f
C13213 a_33496_n8222.t1 VSS 0.021375f
C13214 a_33496_n8222.n2 VSS 0.025404f
C13215 a_33496_n8222.t13 VSS 0.076349f
C13216 a_33496_n8222.t14 VSS 0.04632f
C13217 a_33496_n8222.n3 VSS 0.111235f
C13218 a_33496_n8222.t20 VSS 0.076349f
C13219 a_33496_n8222.t12 VSS 0.04632f
C13220 a_33496_n8222.n4 VSS 0.114323f
C13221 a_33496_n8222.t11 VSS 0.076349f
C13222 a_33496_n8222.t19 VSS 0.04632f
C13223 a_33496_n8222.n5 VSS 0.111235f
C13224 a_33496_n8222.t21 VSS 0.076349f
C13225 a_33496_n8222.t22 VSS 0.04632f
C13226 a_33496_n8222.n6 VSS -0.029833f
C13227 a_33496_n8222.t18 VSS 0.076349f
C13228 a_33496_n8222.t8 VSS 0.04632f
C13229 a_33496_n8222.n7 VSS 0.126528f
C13230 a_33496_n8222.t9 VSS 0.076349f
C13231 a_33496_n8222.t10 VSS 0.04632f
C13232 a_33496_n8222.n8 VSS 0.126528f
C13233 a_33496_n8222.t16 VSS 0.076349f
C13234 a_33496_n8222.t7 VSS 0.04632f
C13235 a_33496_n8222.n9 VSS 0.126528f
C13236 a_33496_n8222.t15 VSS 0.076349f
C13237 a_33496_n8222.t17 VSS 0.04632f
C13238 a_33496_n8222.n10 VSS 0.12344f
C13239 a_33496_n8222.n11 VSS 0.074228f
C13240 a_33496_n8222.n12 VSS 0.058485f
C13241 a_33496_n8222.t6 VSS 0.024116f
C13242 a_21772_n11428.n0 VSS 0.38344f
C13243 a_21772_n11428.t4 VSS 0.019652f
C13244 a_21772_n11428.t6 VSS 0.019652f
C13245 a_21772_n11428.t5 VSS 0.027211f
C13246 a_21772_n11428.n1 VSS 0.047321f
C13247 a_21772_n11428.t3 VSS 0.013209f
C13248 a_21772_n11428.t2 VSS 0.013209f
C13249 a_21772_n11428.n2 VSS 0.026494f
C13250 a_21772_n11428.t1 VSS 0.013209f
C13251 a_21772_n11428.t0 VSS 0.013209f
C13252 a_21772_n11428.n3 VSS 0.031906f
C13253 a_21772_n11428.t22 VSS 0.058056f
C13254 a_21772_n11428.t15 VSS 0.055202f
C13255 a_21772_n11428.n4 VSS 0.090091f
C13256 a_21772_n11428.t18 VSS 0.058056f
C13257 a_21772_n11428.t11 VSS 0.055202f
C13258 a_21772_n11428.n5 VSS 0.090091f
C13259 a_21772_n11428.t21 VSS 0.058056f
C13260 a_21772_n11428.t8 VSS 0.055202f
C13261 a_21772_n11428.n6 VSS -0.035108f
C13262 a_21772_n11428.t23 VSS 0.058056f
C13263 a_21772_n11428.t16 VSS 0.055202f
C13264 a_21772_n11428.n7 VSS 0.101689f
C13265 a_21772_n11428.t19 VSS 0.058056f
C13266 a_21772_n11428.t12 VSS 0.055202f
C13267 a_21772_n11428.n8 VSS 0.101689f
C13268 a_21772_n11428.t14 VSS 0.058056f
C13269 a_21772_n11428.t9 VSS 0.055202f
C13270 a_21772_n11428.n9 VSS 0.101689f
C13271 a_21772_n11428.t17 VSS 0.058056f
C13272 a_21772_n11428.t10 VSS 0.055202f
C13273 a_21772_n11428.n10 VSS 0.101689f
C13274 a_21772_n11428.t20 VSS 0.058056f
C13275 a_21772_n11428.t13 VSS 0.055202f
C13276 a_21772_n11428.n11 VSS 0.146163f
C13277 a_21772_n11428.n12 VSS 0.060222f
C13278 a_21772_n11428.t7 VSS 0.027211f
C13279 OUT[1].t5 VSS 0.014418f
C13280 OUT[1].t2 VSS 0.014418f
C13281 OUT[1].n0 VSS 0.028936f
C13282 OUT[1].t1 VSS 0.014418f
C13283 OUT[1].t7 VSS 0.014418f
C13284 OUT[1].n1 VSS 0.028936f
C13285 OUT[1].t0 VSS 0.014418f
C13286 OUT[1].t4 VSS 0.014418f
C13287 OUT[1].n2 VSS 0.034676f
C13288 OUT[1].n3 VSS 0.158367f
C13289 OUT[1].t8 VSS 0.029702f
C13290 OUT[1].t13 VSS 0.021451f
C13291 OUT[1].n4 VSS 0.051794f
C13292 OUT[1].t9 VSS 0.021451f
C13293 OUT[1].t14 VSS 0.029702f
C13294 OUT[1].n5 VSS 0.064598f
C13295 OUT[1].n6 VSS 0.162514f
C13296 OUT[1].t12 VSS 0.029702f
C13297 OUT[1].t10 VSS 0.021451f
C13298 OUT[1].n7 VSS 0.051794f
C13299 OUT[1].t11 VSS 0.029702f
C13300 OUT[1].t15 VSS 0.021451f
C13301 OUT[1].n8 VSS 0.06552f
C13302 OUT[1].n9 VSS 0.165704f
C13303 OUT[1].n10 VSS 0.127355f
C13304 OUT[1].n11 VSS 0.127355f
C13305 OUT[1].n12 VSS 0.090841f
C13306 OUT[1].t6 VSS 0.014418f
C13307 OUT[1].t3 VSS 0.014418f
C13308 OUT[1].n13 VSS 0.028836f
C13309 OUT[1].n14 VSS 0.371073f
C13310 a_33216_1944.n0 VSS 0.383348f
C13311 a_33216_1944.t5 VSS 0.019652f
C13312 a_33216_1944.t6 VSS 0.027211f
C13313 a_33216_1944.t4 VSS 0.019652f
C13314 a_33216_1944.n1 VSS 0.047321f
C13315 a_33216_1944.t3 VSS 0.013209f
C13316 a_33216_1944.t1 VSS 0.013209f
C13317 a_33216_1944.n2 VSS 0.026494f
C13318 a_33216_1944.t0 VSS 0.013209f
C13319 a_33216_1944.t2 VSS 0.013209f
C13320 a_33216_1944.n3 VSS 0.031906f
C13321 a_33216_1944.t20 VSS 0.055202f
C13322 a_33216_1944.t13 VSS 0.058056f
C13323 a_33216_1944.n4 VSS 0.090091f
C13324 a_33216_1944.t16 VSS 0.055202f
C13325 a_33216_1944.t8 VSS 0.058056f
C13326 a_33216_1944.n5 VSS -0.035108f
C13327 a_33216_1944.t19 VSS 0.055202f
C13328 a_33216_1944.t12 VSS 0.058056f
C13329 a_33216_1944.n6 VSS 0.101689f
C13330 a_33216_1944.t10 VSS 0.055202f
C13331 a_33216_1944.t21 VSS 0.058056f
C13332 a_33216_1944.n7 VSS 0.101689f
C13333 a_33216_1944.t15 VSS 0.055202f
C13334 a_33216_1944.t23 VSS 0.058056f
C13335 a_33216_1944.n8 VSS 0.101689f
C13336 a_33216_1944.t18 VSS 0.055202f
C13337 a_33216_1944.t11 VSS 0.058056f
C13338 a_33216_1944.n9 VSS 0.101689f
C13339 a_33216_1944.t17 VSS 0.055202f
C13340 a_33216_1944.t9 VSS 0.058056f
C13341 a_33216_1944.n10 VSS 0.090091f
C13342 a_33216_1944.t14 VSS 0.055202f
C13343 a_33216_1944.t22 VSS 0.058056f
C13344 a_33216_1944.n11 VSS 0.146257f
C13345 a_33216_1944.n12 VSS 0.060222f
C13346 a_33216_1944.t7 VSS 0.027211f
C13347 a_3935_4156.n0 VSS 0.083919f
C13348 a_3935_4156.n1 VSS 0.086778f
C13349 a_3935_4156.n2 VSS 0.260894f
C13350 a_3935_4156.n3 VSS 1.10322f
C13351 a_3935_4156.t0 VSS 0.086392f
C13352 a_3935_4156.t2 VSS 0.065123f
C13353 a_3935_4156.t13 VSS 0.022527f
C13354 a_3935_4156.t14 VSS 0.022462f
C13355 a_3935_4156.t4 VSS 0.022462f
C13356 a_3935_4156.t5 VSS 0.022462f
C13357 a_3935_4156.t7 VSS 0.022462f
C13358 a_3935_4156.t11 VSS 0.022462f
C13359 a_3935_4156.t6 VSS 0.022462f
C13360 a_3935_4156.t10 VSS 0.022462f
C13361 a_3935_4156.t12 VSS 0.022462f
C13362 a_3935_4156.t3 VSS 0.022462f
C13363 a_3935_4156.t8 VSS 0.028416f
C13364 a_3935_4156.t9 VSS 0.042963f
C13365 a_3935_4156.n4 VSS 0.155027f
C13366 a_3935_4156.n5 VSS 0.290234f
C13367 a_3935_4156.t1 VSS 0.072354f
C13368 a_13501_n17172.n0 VSS 2.0189f
C13369 a_13501_n17172.n1 VSS 3.79312f
C13370 a_13501_n17172.t17 VSS 0.33153f
C13371 a_13501_n17172.t9 VSS 0.321965f
C13372 a_13501_n17172.t7 VSS 0.041646f
C13373 a_13501_n17172.t1 VSS 0.041646f
C13374 a_13501_n17172.n2 VSS 0.229216f
C13375 a_13501_n17172.t15 VSS 0.041646f
C13376 a_13501_n17172.t19 VSS 0.041646f
C13377 a_13501_n17172.n3 VSS 0.223712f
C13378 a_13501_n17172.t4 VSS 0.041646f
C13379 a_13501_n17172.t8 VSS 0.041646f
C13380 a_13501_n17172.n4 VSS 0.228449f
C13381 a_13501_n17172.t12 VSS 0.041646f
C13382 a_13501_n17172.t16 VSS 0.041646f
C13383 a_13501_n17172.n5 VSS 0.22515f
C13384 a_13501_n17172.t10 VSS 0.041646f
C13385 a_13501_n17172.t13 VSS 0.041646f
C13386 a_13501_n17172.n6 VSS 0.22515f
C13387 a_13501_n17172.t2 VSS 0.041646f
C13388 a_13501_n17172.t5 VSS 0.041646f
C13389 a_13501_n17172.n7 VSS 0.227874f
C13390 a_13501_n17172.t3 VSS 0.041646f
C13391 a_13501_n17172.t6 VSS 0.041646f
C13392 a_13501_n17172.n8 VSS 0.228065f
C13393 a_13501_n17172.t11 VSS 0.041646f
C13394 a_13501_n17172.t14 VSS 0.041646f
C13395 a_13501_n17172.n9 VSS 0.22387f
C13396 a_13501_n17172.t0 VSS 0.325425f
C13397 a_13501_n17172.t18 VSS 0.33124f
C13398 a_21996_332.n0 VSS 1.30554f
C13399 a_21996_332.t1 VSS 0.024343f
C13400 a_21996_332.t0 VSS 0.015657f
C13401 a_21996_332.t3 VSS 0.020404f
C13402 a_21996_332.t2 VSS 0.0245f
C13403 a_21996_332.n1 VSS 1.00956f
C13404 a_29076_n8292.t2 VSS 0.048847f
C13405 a_29076_n8292.t3 VSS 0.043605f
C13406 a_29076_n8292.t0 VSS 0.046911f
C13407 a_29076_n8292.t1 VSS 0.043605f
C13408 a_29076_n8292.n0 VSS 0.243969f
C13409 a_29076_n8292.t7 VSS 0.041313f
C13410 a_29076_n8292.t9 VSS 0.037565f
C13411 a_29076_n8292.n1 VSS 0.047532f
C13412 a_29076_n8292.t10 VSS 0.029768f
C13413 a_29076_n8292.t4 VSS 0.031074f
C13414 a_29076_n8292.n2 VSS 0.069375f
C13415 a_29076_n8292.n3 VSS 0.240745f
C13416 a_29076_n8292.t6 VSS 0.039721f
C13417 a_29076_n8292.t8 VSS 0.036011f
C13418 a_29076_n8292.n4 VSS 0.166583f
C13419 a_29076_n8292.n5 VSS 0.808783f
C13420 a_29076_n8292.t11 VSS 0.046108f
C13421 a_29076_n8292.t5 VSS 0.030265f
C13422 a_29076_n8292.n6 VSS 0.191515f
C13423 a_29076_n8292.n7 VSS 0.556702f
C13424 a_34708_n5896.n0 VSS 0.297367f
C13425 a_34708_n5896.n1 VSS 0.551684f
C13426 a_34708_n5896.n2 VSS 0.207454f
C13427 a_34708_n5896.t9 VSS 0.043182f
C13428 a_34708_n5896.t11 VSS 0.043182f
C13429 a_34708_n5896.t14 VSS 0.043182f
C13430 a_34708_n5896.n3 VSS 0.107923f
C13431 a_34708_n5896.t12 VSS 0.043182f
C13432 a_34708_n5896.t10 VSS 0.043182f
C13433 a_34708_n5896.n4 VSS 0.087445f
C13434 a_34708_n5896.t13 VSS 0.043182f
C13435 a_34708_n5896.t8 VSS 0.043182f
C13436 a_34708_n5896.n5 VSS 0.107923f
C13437 a_34708_n5896.t1 VSS 0.010992f
C13438 a_34708_n5896.t7 VSS 0.010992f
C13439 a_34708_n5896.n6 VSS 0.022326f
C13440 a_34708_n5896.t0 VSS 0.010992f
C13441 a_34708_n5896.t6 VSS 0.010992f
C13442 a_34708_n5896.n7 VSS 0.031493f
C13443 a_34708_n5896.t2 VSS 0.010992f
C13444 a_34708_n5896.t5 VSS 0.010992f
C13445 a_34708_n5896.n8 VSS 0.022326f
C13446 a_34708_n5896.t3 VSS 0.010992f
C13447 a_34708_n5896.t4 VSS 0.010992f
C13448 a_34708_n5896.n9 VSS 0.031493f
C13449 a_34708_n5896.t27 VSS 0.124345f
C13450 a_34708_n5896.t20 VSS 0.081985f
C13451 a_34708_n5896.t26 VSS 0.046013f
C13452 a_34708_n5896.n10 VSS 0.219353f
C13453 a_34708_n5896.t29 VSS 0.081985f
C13454 a_34708_n5896.t21 VSS 0.046013f
C13455 a_34708_n5896.n11 VSS 0.141711f
C13456 a_34708_n5896.t25 VSS 0.081985f
C13457 a_34708_n5896.t18 VSS 0.046013f
C13458 a_34708_n5896.n12 VSS 0.14879f
C13459 a_34708_n5896.n13 VSS 0.276066f
C13460 a_34708_n5896.t16 VSS 0.081985f
C13461 a_34708_n5896.t24 VSS 0.046013f
C13462 a_34708_n5896.n14 VSS 0.141711f
C13463 a_34708_n5896.t19 VSS 0.081985f
C13464 a_34708_n5896.t22 VSS 0.046013f
C13465 a_34708_n5896.n15 VSS 0.14879f
C13466 a_34708_n5896.t17 VSS 0.124345f
C13467 a_34708_n5896.t28 VSS 0.081985f
C13468 a_34708_n5896.t23 VSS 0.046013f
C13469 a_34708_n5896.n16 VSS 0.219353f
C13470 a_34708_n5896.n17 VSS 0.382946f
C13471 a_34708_n5896.n18 VSS 0.816328f
C13472 a_34708_n5896.n19 VSS 0.087445f
C13473 a_34708_n5896.t15 VSS 0.043182f
C13474 a_33776_n5896.n0 VSS 0.466769f
C13475 a_33776_n5896.t4 VSS 0.024116f
C13476 a_33776_n5896.t5 VSS 0.024116f
C13477 a_33776_n5896.t3 VSS 0.024116f
C13478 a_33776_n5896.n1 VSS 0.04873f
C13479 a_33776_n5896.t0 VSS 0.021374f
C13480 a_33776_n5896.n2 VSS 0.025404f
C13481 a_33776_n5896.t14 VSS 0.04632f
C13482 a_33776_n5896.t17 VSS 0.076349f
C13483 a_33776_n5896.n3 VSS 0.111235f
C13484 a_33776_n5896.t13 VSS 0.04632f
C13485 a_33776_n5896.t9 VSS 0.076349f
C13486 a_33776_n5896.n4 VSS -0.029833f
C13487 a_33776_n5896.t16 VSS 0.04632f
C13488 a_33776_n5896.t19 VSS 0.076349f
C13489 a_33776_n5896.n5 VSS 0.126528f
C13490 a_33776_n5896.t12 VSS 0.04632f
C13491 a_33776_n5896.t8 VSS 0.076349f
C13492 a_33776_n5896.n6 VSS 0.126528f
C13493 a_33776_n5896.t21 VSS 0.04632f
C13494 a_33776_n5896.t15 VSS 0.076349f
C13495 a_33776_n5896.n7 VSS 0.126528f
C13496 a_33776_n5896.t7 VSS 0.04632f
C13497 a_33776_n5896.t18 VSS 0.076349f
C13498 a_33776_n5896.n8 VSS 0.12344f
C13499 a_33776_n5896.t10 VSS 0.04632f
C13500 a_33776_n5896.t20 VSS 0.076349f
C13501 a_33776_n5896.n9 VSS 0.111235f
C13502 a_33776_n5896.t22 VSS 0.04632f
C13503 a_33776_n5896.t11 VSS 0.076349f
C13504 a_33776_n5896.n10 VSS 0.114323f
C13505 a_33776_n5896.n11 VSS 0.074228f
C13506 a_33776_n5896.n12 VSS 0.058485f
C13507 a_33776_n5896.t6 VSS 0.024116f
C13508 a_13501_n14494.n0 VSS 2.0189f
C13509 a_13501_n14494.n1 VSS 3.79312f
C13510 a_13501_n14494.t11 VSS 0.041646f
C13511 a_13501_n14494.t15 VSS 0.33153f
C13512 a_13501_n14494.t3 VSS 0.321965f
C13513 a_13501_n14494.t5 VSS 0.041646f
C13514 a_13501_n14494.t1 VSS 0.041646f
C13515 a_13501_n14494.n2 VSS 0.229216f
C13516 a_13501_n14494.t13 VSS 0.041646f
C13517 a_13501_n14494.t17 VSS 0.041646f
C13518 a_13501_n14494.n3 VSS 0.223712f
C13519 a_13501_n14494.t8 VSS 0.041646f
C13520 a_13501_n14494.t4 VSS 0.041646f
C13521 a_13501_n14494.n4 VSS 0.228449f
C13522 a_13501_n14494.t10 VSS 0.041646f
C13523 a_13501_n14494.t14 VSS 0.041646f
C13524 a_13501_n14494.n5 VSS 0.22515f
C13525 a_13501_n14494.t16 VSS 0.33124f
C13526 a_13501_n14494.t2 VSS 0.325425f
C13527 a_13501_n14494.t19 VSS 0.041646f
C13528 a_13501_n14494.t12 VSS 0.041646f
C13529 a_13501_n14494.n6 VSS 0.22387f
C13530 a_13501_n14494.t9 VSS 0.041646f
C13531 a_13501_n14494.t6 VSS 0.041646f
C13532 a_13501_n14494.n7 VSS 0.228065f
C13533 a_13501_n14494.t0 VSS 0.041646f
C13534 a_13501_n14494.t7 VSS 0.041646f
C13535 a_13501_n14494.n8 VSS 0.227874f
C13536 a_13501_n14494.n9 VSS 0.22515f
C13537 a_13501_n14494.t18 VSS 0.041646f
C13538 a_4001_4292.n0 VSS 0.101735f
C13539 a_4001_4292.n1 VSS 0.105241f
C13540 a_4001_4292.n2 VSS 0.158385f
C13541 a_4001_4292.t0 VSS 0.071534f
C13542 a_4001_4292.t4 VSS 0.026854f
C13543 a_4001_4292.t5 VSS 0.026778f
C13544 a_4001_4292.t3 VSS 0.026778f
C13545 a_4001_4292.t7 VSS 0.026778f
C13546 a_4001_4292.t8 VSS 0.026778f
C13547 a_4001_4292.t9 VSS 0.026778f
C13548 a_4001_4292.t10 VSS 0.026778f
C13549 a_4001_4292.t13 VSS 0.026778f
C13550 a_4001_4292.t11 VSS 0.026778f
C13551 a_4001_4292.t12 VSS 0.026778f
C13552 a_4001_4292.t6 VSS 0.049784f
C13553 a_4001_4292.t14 VSS 0.033875f
C13554 a_4001_4292.n3 VSS 0.961573f
C13555 a_4001_4292.n4 VSS 0.18446f
C13556 a_4001_4292.t2 VSS 0.099908f
C13557 a_4001_4292.n5 VSS 0.378197f
C13558 a_4001_4292.t1 VSS 0.087456f
C13559 a_25020_n8200.t1 VSS 0.143937f
C13560 a_25020_n8200.n0 VSS 1.54412f
C13561 a_25020_n8200.t0 VSS 0.023601f
C13562 a_25020_n8200.t4 VSS 0.018085f
C13563 a_25020_n8200.t6 VSS 0.036603f
C13564 a_25020_n8200.n1 VSS 0.322998f
C13565 a_25020_n8200.t7 VSS 0.037747f
C13566 a_25020_n8200.t3 VSS 0.020529f
C13567 a_25020_n8200.n2 VSS 0.088566f
C13568 a_25020_n8200.t5 VSS 0.029099f
C13569 a_25020_n8200.t2 VSS 0.01853f
C13570 a_25020_n8200.n3 VSS 0.216185f
C13571 a_13623_n20230.n0 VSS 4.01842f
C13572 a_13623_n20230.n1 VSS 5.46815f
C13573 a_13623_n20230.n2 VSS 0.476923f
C13574 a_13623_n20230.n3 VSS 0.084936f
C13575 a_13623_n20230.n4 VSS 0.32079f
C13576 a_13623_n20230.t9 VSS 0.016211f
C13577 a_13623_n20230.t12 VSS 0.011708f
C13578 a_13623_n20230.t14 VSS 0.016211f
C13579 a_13623_n20230.n5 VSS 0.028269f
C13580 a_13623_n20230.t13 VSS 0.016211f
C13581 a_13623_n20230.t11 VSS 0.011708f
C13582 a_13623_n20230.n6 VSS 0.035257f
C13583 a_13623_n20230.n7 VSS 0.015793f
C13584 a_13623_n20230.n8 VSS 0.018926f
C13585 a_13623_n20230.n9 VSS 0.015793f
C13586 a_13623_n20230.n10 VSS 0.018988f
C13587 a_13623_n20230.t8 VSS 0.011708f
C13588 a_13623_n20230.t10 VSS 0.016211f
C13589 a_13623_n20230.n11 VSS 0.028269f
C13590 a_13623_n20230.t29 VSS 0.045486f
C13591 a_13623_n20230.t26 VSS 0.04566f
C13592 a_13623_n20230.t16 VSS 0.045486f
C13593 a_13623_n20230.t36 VSS 0.045486f
C13594 a_13623_n20230.t24 VSS 0.045486f
C13595 a_13623_n20230.t45 VSS 0.045486f
C13596 a_13623_n20230.t23 VSS 0.045486f
C13597 a_13623_n20230.t38 VSS 0.045486f
C13598 a_13623_n20230.t30 VSS 0.045486f
C13599 a_13623_n20230.t17 VSS 0.045486f
C13600 a_13623_n20230.t33 VSS 0.045745f
C13601 a_13623_n20230.t42 VSS 0.045651f
C13602 a_13623_n20230.t25 VSS 0.045486f
C13603 a_13623_n20230.t34 VSS 0.045486f
C13604 a_13623_n20230.t28 VSS 0.045486f
C13605 a_13623_n20230.t39 VSS 0.045486f
C13606 a_13623_n20230.t20 VSS 0.045486f
C13607 a_13623_n20230.t31 VSS 0.045486f
C13608 a_13623_n20230.t41 VSS 0.045486f
C13609 a_13623_n20230.t22 VSS 0.045486f
C13610 a_13623_n20230.t18 VSS 0.045486f
C13611 a_13623_n20230.t37 VSS 0.045508f
C13612 a_13623_n20230.t44 VSS 0.04566f
C13613 a_13623_n20230.t27 VSS 0.04566f
C13614 a_13623_n20230.t35 VSS 0.04566f
C13615 a_13623_n20230.t19 VSS 0.04566f
C13616 a_13623_n20230.t40 VSS 0.04566f
C13617 a_13623_n20230.t21 VSS 0.04566f
C13618 a_13623_n20230.t32 VSS 0.04566f
C13619 a_13623_n20230.t43 VSS 0.04566f
C13620 a_13623_n20230.n12 VSS 0.028269f
C13621 a_13623_n20230.t15 VSS 0.011708f
C13622 a_21772_n3588.n0 VSS 0.61362f
C13623 a_21772_n3588.t0 VSS 0.055212f
C13624 a_21772_n3588.t2 VSS 0.060859f
C13625 a_21772_n3588.t1 VSS 0.067887f
C13626 a_21772_n3588.t3 VSS 0.081141f
C13627 a_21772_n3588.t9 VSS 0.06058f
C13628 a_21772_n3588.t7 VSS 0.057602f
C13629 a_21772_n3588.n1 VSS 0.094008f
C13630 a_21772_n3588.t13 VSS 0.06058f
C13631 a_21772_n3588.t12 VSS 0.057602f
C13632 a_21772_n3588.n2 VSS 0.094008f
C13633 a_21772_n3588.t19 VSS 0.06058f
C13634 a_21772_n3588.t14 VSS 0.057602f
C13635 a_21772_n3588.n3 VSS -0.036634f
C13636 a_21772_n3588.t16 VSS 0.06058f
C13637 a_21772_n3588.t15 VSS 0.057602f
C13638 a_21772_n3588.n4 VSS 0.106111f
C13639 a_21772_n3588.t4 VSS 0.06058f
C13640 a_21772_n3588.t17 VSS 0.057602f
C13641 a_21772_n3588.n5 VSS 0.106111f
C13642 a_21772_n3588.t6 VSS 0.06058f
C13643 a_21772_n3588.t5 VSS 0.057602f
C13644 a_21772_n3588.n6 VSS 0.106111f
C13645 a_21772_n3588.t10 VSS 0.06058f
C13646 a_21772_n3588.t18 VSS 0.057602f
C13647 a_21772_n3588.n7 VSS 0.106111f
C13648 a_21772_n3588.t11 VSS 0.06058f
C13649 a_21772_n3588.t8 VSS 0.057602f
C13650 a_29920_n3900.t0 VSS 0.094024f
C13651 a_29920_n3900.n0 VSS 1.74669f
C13652 a_29920_n3900.n1 VSS 0.142069f
C13653 a_29920_n3900.t1 VSS 0.143502f
C13654 a_29920_n3900.n3 VSS 0.583578f
C13655 a_29920_n3900.n4 VSS 0.154876f
C13656 a_29920_n3900.t13 VSS 0.100875f
C13657 a_29920_n3900.t18 VSS 0.049841f
C13658 a_29920_n3900.n5 VSS 0.510043f
C13659 a_29920_n3900.t2 VSS 0.06147f
C13660 a_29920_n3900.t17 VSS 0.098464f
C13661 a_29920_n3900.n6 VSS 0.142079f
C13662 a_29920_n3900.t7 VSS 0.06147f
C13663 a_29920_n3900.t14 VSS 0.098464f
C13664 a_29920_n3900.n7 VSS 0.142079f
C13665 a_29920_n3900.t23 VSS 0.06147f
C13666 a_29920_n3900.t10 VSS 0.098464f
C13667 a_29920_n3900.n8 VSS 0.5173f
C13668 a_29920_n3900.t16 VSS 0.081325f
C13669 a_29920_n3900.t21 VSS 0.104552f
C13670 a_29920_n3900.n9 VSS 0.932052f
C13671 a_29920_n3900.t20 VSS 0.088003f
C13672 a_29920_n3900.t9 VSS 0.101298f
C13673 a_29920_n3900.n10 VSS 0.135857f
C13674 a_29920_n3900.t12 VSS 0.088003f
C13675 a_29920_n3900.t15 VSS 0.087916f
C13676 a_29920_n3900.t8 VSS 0.093624f
C13677 a_29920_n3900.t5 VSS 0.095207f
C13678 a_29920_n3900.t11 VSS 0.088003f
C13679 a_29920_n3900.t3 VSS 0.101298f
C13680 a_29920_n3900.n11 VSS 0.123553f
C13681 a_29920_n3900.n12 VSS 1.02105f
C13682 a_29920_n3900.t19 VSS 0.078478f
C13683 a_29920_n3900.t22 VSS 0.104027f
C13684 a_29920_n3900.n13 VSS 0.132524f
C13685 a_29920_n3900.t4 VSS 0.104733f
C13686 a_29920_n3900.t6 VSS 0.08091f
C13687 a_29920_n3900.n14 VSS 0.130753f
C13688 a_29920_n3900.n15 VSS 0.214897f
C13689 a_29920_n3900.n16 VSS 0.392087f
C13690 a_29920_n3900.n17 VSS 0.313085f
C13691 a_23072_n13432.n0 VSS 0.254851f
C13692 a_23072_n13432.n1 VSS 0.459823f
C13693 a_23072_n13432.t1 VSS 0.023535f
C13694 a_23072_n13432.t3 VSS 0.028405f
C13695 a_23072_n13432.t2 VSS 0.028405f
C13696 a_23072_n13432.t4 VSS 0.023535f
C13697 a_23072_n13432.n2 VSS 0.989895f
C13698 a_23072_n13432.n3 VSS 0.064446f
C13699 a_23072_n13432.n4 VSS 0.64295f
C13700 a_23072_n13432.n5 VSS 0.739157f
C13701 a_23072_n13432.n6 VSS 0.492356f
C13702 a_23072_n13432.n7 VSS 0.629282f
C13703 a_23072_n13432.n8 VSS 0.686817f
C13704 a_23072_n13432.t0 VSS 0.092318f
C13705 a_23072_n13432.n9 VSS 0.68981f
C13706 a_23072_n13432.n10 VSS 0.064446f
C13707 a_23072_n13432.n11 VSS 0.318576f
C13708 a_23072_n13432.n12 VSS 0.356255f
C13709 a_23072_n13432.t6 VSS 0.063302f
C13710 a_23072_n13432.t5 VSS 0.062343f
C13711 a_23072_n13432.t7 VSS 0.072557f
C13712 a_23072_n13432.t44 VSS 0.023911f
C13713 a_23072_n13432.t72 VSS 0.021432f
C13714 a_23072_n13432.n13 VSS 0.131451f
C13715 a_23072_n13432.t64 VSS 0.023459f
C13716 a_23072_n13432.t27 VSS 0.021438f
C13717 a_23072_n13432.n14 VSS 0.252379f
C13718 a_23072_n13432.t28 VSS 0.023911f
C13719 a_23072_n13432.t33 VSS 0.021432f
C13720 a_23072_n13432.n15 VSS 0.059662f
C13721 a_23072_n13432.n16 VSS 1.13242f
C13722 a_23072_n13432.t76 VSS 0.021438f
C13723 a_23072_n13432.t80 VSS 0.023459f
C13724 a_23072_n13432.t102 VSS 0.065015f
C13725 a_23072_n13432.t40 VSS 0.062077f
C13726 a_23072_n13432.t66 VSS 0.182584f
C13727 a_23072_n13432.t45 VSS 0.137161f
C13728 a_23072_n13432.n17 VSS 0.149679f
C13729 a_23072_n13432.t99 VSS 0.062077f
C13730 a_23072_n13432.t21 VSS 0.182584f
C13731 a_23072_n13432.t68 VSS 0.137161f
C13732 a_23072_n13432.t61 VSS 0.065015f
C13733 a_23072_n13432.n18 VSS 0.087914f
C13734 a_23072_n13432.t17 VSS 0.021438f
C13735 a_23072_n13432.t8 VSS 0.023459f
C13736 a_23072_n13432.t55 VSS 0.062077f
C13737 a_23072_n13432.t79 VSS 0.182584f
C13738 a_23072_n13432.t59 VSS 0.137161f
C13739 a_23072_n13432.t35 VSS 0.065015f
C13740 a_23072_n13432.n19 VSS 0.058412f
C13741 a_23072_n13432.t20 VSS 0.022872f
C13742 a_23072_n13432.t92 VSS 0.021666f
C13743 a_23072_n13432.n20 VSS 0.116905f
C13744 a_23072_n13432.t51 VSS 0.0219f
C13745 a_23072_n13432.t16 VSS 0.022358f
C13746 a_23072_n13432.t22 VSS 0.0219f
C13747 a_23072_n13432.t89 VSS 0.022358f
C13748 a_23072_n13432.n21 VSS 0.237092f
C13749 a_23072_n13432.n22 VSS 0.347596f
C13750 a_23072_n13432.t100 VSS 0.021438f
C13751 a_23072_n13432.t74 VSS 0.023459f
C13752 a_23072_n13432.t56 VSS 0.023459f
C13753 a_23072_n13432.t15 VSS 0.021438f
C13754 a_23072_n13432.n23 VSS 0.101693f
C13755 a_23072_n13432.t54 VSS 0.0219f
C13756 a_23072_n13432.t52 VSS 0.022358f
C13757 a_23072_n13432.n24 VSS 0.077606f
C13758 a_23072_n13432.t77 VSS 0.065015f
C13759 a_23072_n13432.t29 VSS 0.062077f
C13760 a_23072_n13432.t23 VSS 0.182584f
C13761 a_23072_n13432.t85 VSS 0.137161f
C13762 a_23072_n13432.n25 VSS 0.333893f
C13763 a_23072_n13432.t26 VSS 0.062077f
C13764 a_23072_n13432.t94 VSS 0.182584f
C13765 a_23072_n13432.t30 VSS 0.137161f
C13766 a_23072_n13432.t48 VSS 0.065015f
C13767 a_23072_n13432.n26 VSS 0.089491f
C13768 a_23072_n13432.n27 VSS 0.793897f
C13769 a_23072_n13432.t71 VSS 0.023911f
C13770 a_23072_n13432.t60 VSS 0.021432f
C13771 a_23072_n13432.n28 VSS 0.201367f
C13772 a_23072_n13432.t95 VSS 0.062077f
C13773 a_23072_n13432.t93 VSS 0.182584f
C13774 a_23072_n13432.t10 VSS 0.137161f
C13775 a_23072_n13432.t57 VSS 0.065015f
C13776 a_23072_n13432.n29 VSS 0.110135f
C13777 a_23072_n13432.n30 VSS 0.863369f
C13778 a_23072_n13432.t42 VSS 0.021666f
C13779 a_23072_n13432.t87 VSS 0.022872f
C13780 a_23072_n13432.n31 VSS 0.072408f
C13781 a_23072_n13432.n32 VSS 0.568567f
C13782 a_23072_n13432.t18 VSS 0.062077f
C13783 a_23072_n13432.t103 VSS 0.182584f
C13784 a_23072_n13432.t91 VSS 0.137161f
C13785 a_23072_n13432.t69 VSS 0.065015f
C13786 a_23072_n13432.n33 VSS 0.1168f
C13787 a_23072_n13432.n34 VSS 0.431159f
C13788 a_23072_n13432.t86 VSS 0.030641f
C13789 a_23072_n13432.t43 VSS 0.067543f
C13790 a_23072_n13432.t53 VSS 0.1561f
C13791 a_23072_n13432.t101 VSS 0.120857f
C13792 a_23072_n13432.n35 VSS 0.068357f
C13793 a_23072_n13432.t82 VSS 0.062077f
C13794 a_23072_n13432.t65 VSS 0.182584f
C13795 a_23072_n13432.t84 VSS 0.137161f
C13796 a_23072_n13432.t14 VSS 0.065015f
C13797 a_23072_n13432.n36 VSS 0.088414f
C13798 a_23072_n13432.t25 VSS 0.062077f
C13799 a_23072_n13432.t98 VSS 0.182584f
C13800 a_23072_n13432.t38 VSS 0.137161f
C13801 a_23072_n13432.t73 VSS 0.065015f
C13802 a_23072_n13432.n37 VSS 0.058769f
C13803 a_23072_n13432.n38 VSS 0.500677f
C13804 a_23072_n13432.t24 VSS 0.062077f
C13805 a_23072_n13432.t97 VSS 0.182584f
C13806 a_23072_n13432.t37 VSS 0.137161f
C13807 a_23072_n13432.t62 VSS 0.065015f
C13808 a_23072_n13432.n39 VSS 0.087914f
C13809 a_23072_n13432.n40 VSS 0.295055f
C13810 a_23072_n13432.t46 VSS 0.023459f
C13811 a_23072_n13432.t32 VSS 0.021438f
C13812 a_23072_n13432.n41 VSS 0.078723f
C13813 a_23072_n13432.t96 VSS 0.023911f
C13814 a_23072_n13432.t88 VSS 0.021432f
C13815 a_23072_n13432.n42 VSS 0.142063f
C13816 a_23072_n13432.t70 VSS 0.062077f
C13817 a_23072_n13432.t9 VSS 0.182584f
C13818 a_23072_n13432.t49 VSS 0.137161f
C13819 a_23072_n13432.t50 VSS 0.065015f
C13820 a_23072_n13432.n43 VSS 0.123826f
C13821 a_23072_n13432.t12 VSS 0.062077f
C13822 a_23072_n13432.t58 VSS 0.182584f
C13823 a_23072_n13432.t13 VSS 0.137161f
C13824 a_23072_n13432.t34 VSS 0.065015f
C13825 a_23072_n13432.n44 VSS 0.087914f
C13826 a_23072_n13432.t47 VSS 0.062077f
C13827 a_23072_n13432.t75 VSS 0.182584f
C13828 a_23072_n13432.t11 VSS 0.137161f
C13829 a_23072_n13432.t19 VSS 0.065015f
C13830 a_23072_n13432.n45 VSS 0.090763f
C13831 a_23072_n13432.n46 VSS 0.302543f
C13832 a_23072_n13432.t41 VSS 0.065015f
C13833 a_23072_n13432.t31 VSS 0.062077f
C13834 a_23072_n13432.t39 VSS 0.182584f
C13835 a_23072_n13432.t67 VSS 0.137161f
C13836 a_23072_n13432.n47 VSS 0.128876f
C13837 a_23072_n13432.n48 VSS 0.509362f
C13838 a_23072_n13432.n49 VSS 0.354333f
C13839 a_23072_n13432.t81 VSS 0.065015f
C13840 a_23072_n13432.t36 VSS 0.062077f
C13841 a_23072_n13432.t63 VSS 0.182584f
C13842 a_23072_n13432.t83 VSS 0.137161f
C13843 a_23072_n13432.n50 VSS 0.110135f
C13844 a_23072_n13432.t90 VSS 0.023911f
C13845 a_23072_n13432.t78 VSS 0.021432f
C13846 a_23072_n13432.n51 VSS 0.059662f
C13847 a_11023_n9518.n0 VSS 0.016468f
C13848 a_11023_n9518.n1 VSS 0.640198f
C13849 a_11023_n9518.n2 VSS 0.056878f
C13850 a_11023_n9518.n3 VSS 0.016571f
C13851 a_11023_n9518.n4 VSS 0.056671f
C13852 a_11023_n9518.n5 VSS 0.056464f
C13853 a_11023_n9518.n6 VSS 0.056257f
C13854 a_11023_n9518.n7 VSS 0.315152f
C13855 a_11023_n9518.n8 VSS 0.315152f
C13856 a_11023_n9518.n9 VSS 0.315152f
C13857 a_11023_n9518.n10 VSS 0.436195f
C13858 a_11023_n9518.n11 VSS 0.106969f
C13859 a_11023_n9518.n12 VSS 0.052321f
C13860 a_11023_n9518.n13 VSS 0.021957f
C13861 a_11023_n9518.n14 VSS 0.052114f
C13862 a_11023_n9518.n15 VSS 0.021957f
C13863 a_11023_n9518.n16 VSS 0.051907f
C13864 a_11023_n9518.n17 VSS 0.0517f
C13865 a_11023_n9518.t15 VSS 0.0377f
C13866 a_11023_n9518.t14 VSS 0.0377f
C13867 a_11023_n9518.t18 VSS 0.0377f
C13868 a_11023_n9518.n18 VSS 0.196436f
C13869 a_11023_n9518.t16 VSS 0.0377f
C13870 a_11023_n9518.t12 VSS 0.0377f
C13871 a_11023_n9518.n19 VSS 0.181424f
C13872 a_11023_n9518.n20 VSS 0.503298f
C13873 a_11023_n9518.t22 VSS 0.064188f
C13874 a_11023_n9518.n21 VSS 0.144341f
C13875 a_11023_n9518.t34 VSS 0.064062f
C13876 a_11023_n9518.n22 VSS 0.055918f
C13877 a_11023_n9518.t37 VSS 0.064062f
C13878 a_11023_n9518.n23 VSS 0.016571f
C13879 a_11023_n9518.n24 VSS 0.119271f
C13880 a_11023_n9518.n25 VSS 0.021957f
C13881 a_11023_n9518.n26 VSS 0.021957f
C13882 a_11023_n9518.t23 VSS 0.064062f
C13883 a_11023_n9518.t32 VSS 0.064062f
C13884 a_11023_n9518.t27 VSS 0.064062f
C13885 a_11023_n9518.t20 VSS 0.064062f
C13886 a_11023_n9518.t25 VSS 0.06392f
C13887 a_11023_n9518.t31 VSS 0.063818f
C13888 a_11023_n9518.t39 VSS 0.063818f
C13889 a_11023_n9518.t26 VSS 0.063818f
C13890 a_11023_n9518.t33 VSS 0.063818f
C13891 a_11023_n9518.t21 VSS 0.063818f
C13892 a_11023_n9518.t28 VSS 0.063818f
C13893 a_11023_n9518.t24 VSS 0.063818f
C13894 a_11023_n9518.t29 VSS 0.063818f
C13895 a_11023_n9518.t38 VSS 0.063818f
C13896 a_11023_n9518.n27 VSS 0.221496f
C13897 a_11023_n9518.t30 VSS 0.064062f
C13898 a_11023_n9518.n28 VSS 0.071939f
C13899 a_11023_n9518.n29 VSS 0.021957f
C13900 a_11023_n9518.n30 VSS 0.016571f
C13901 a_11023_n9518.t35 VSS 0.064062f
C13902 a_11023_n9518.n31 VSS 0.021957f
C13903 a_11023_n9518.n32 VSS 0.021957f
C13904 a_11023_n9518.n33 VSS 0.016571f
C13905 a_11023_n9518.t36 VSS 0.064062f
C13906 a_11023_n9518.t2 VSS 0.0377f
C13907 a_11023_n9518.t6 VSS 0.0377f
C13908 a_11023_n9518.n34 VSS 0.179009f
C13909 a_11023_n9518.t5 VSS 0.0377f
C13910 a_11023_n9518.t8 VSS 0.0377f
C13911 a_11023_n9518.n35 VSS 0.179009f
C13912 a_11023_n9518.t4 VSS 0.0377f
C13913 a_11023_n9518.t1 VSS 0.0377f
C13914 a_11023_n9518.n36 VSS 0.179009f
C13915 a_11023_n9518.t7 VSS 0.0377f
C13916 a_11023_n9518.t0 VSS 0.0377f
C13917 a_11023_n9518.n37 VSS 0.179009f
C13918 a_11023_n9518.t9 VSS 0.0377f
C13919 a_11023_n9518.t3 VSS 0.0377f
C13920 a_11023_n9518.n38 VSS 0.198821f
C13921 a_11023_n9518.n39 VSS 0.696191f
C13922 a_11023_n9518.n40 VSS 0.29804f
C13923 a_11023_n9518.n41 VSS 0.29804f
C13924 a_11023_n9518.n42 VSS 0.414463f
C13925 a_11023_n9518.n43 VSS 0.718664f
C13926 a_11023_n9518.t13 VSS 0.0377f
C13927 a_11023_n9518.t11 VSS 0.0377f
C13928 a_11023_n9518.n44 VSS 0.181424f
C13929 a_11023_n9518.n45 VSS 0.319464f
C13930 a_11023_n9518.t10 VSS 0.0377f
C13931 a_11023_n9518.t17 VSS 0.0377f
C13932 a_11023_n9518.n46 VSS 0.181424f
C13933 a_11023_n9518.n47 VSS 0.184638f
C13934 a_11023_n9518.n48 VSS 0.184636f
C13935 a_11023_n9518.n49 VSS 0.181426f
C13936 a_11023_n9518.t19 VSS 0.0377f
C13937 a_13623_n4162.n0 VSS 3.83703f
C13938 a_13623_n4162.n1 VSS 0.448485f
C13939 a_13623_n4162.n2 VSS 0.079872f
C13940 a_13623_n4162.n3 VSS 0.350028f
C13941 a_13623_n4162.n4 VSS 0.301662f
C13942 a_13623_n4162.t9 VSS 0.01101f
C13943 a_13623_n4162.t13 VSS 0.01101f
C13944 a_13623_n4162.t12 VSS 0.015244f
C13945 a_13623_n4162.n5 VSS 0.026583f
C13946 a_13623_n4162.t14 VSS 0.015244f
C13947 a_13623_n4162.t8 VSS 0.01101f
C13948 a_13623_n4162.n6 VSS 0.033155f
C13949 a_13623_n4162.n7 VSS 0.014851f
C13950 a_13623_n4162.n8 VSS 0.017797f
C13951 a_13623_n4162.n9 VSS 0.014851f
C13952 a_13623_n4162.n10 VSS 0.017856f
C13953 a_13623_n4162.t21 VSS 0.042774f
C13954 a_13623_n4162.t23 VSS 0.042937f
C13955 a_13623_n4162.t40 VSS 0.042774f
C13956 a_13623_n4162.t44 VSS 0.042937f
C13957 a_13623_n4162.t16 VSS 0.042774f
C13958 a_13623_n4162.t18 VSS 0.042937f
C13959 a_13623_n4162.t29 VSS 0.042774f
C13960 a_13623_n4162.t33 VSS 0.042937f
C13961 a_13623_n4162.t38 VSS 0.042774f
C13962 a_13623_n4162.t42 VSS 0.042937f
C13963 a_13623_n4162.t17 VSS 0.042774f
C13964 a_13623_n4162.t20 VSS 0.042937f
C13965 a_13623_n4162.t32 VSS 0.042774f
C13966 a_13623_n4162.t37 VSS 0.042937f
C13967 a_13623_n4162.t41 VSS 0.042774f
C13968 a_13623_n4162.t45 VSS 0.042937f
C13969 a_13623_n4162.t24 VSS 0.042774f
C13970 a_13623_n4162.t35 VSS 0.043018f
C13971 a_13623_n4162.t22 VSS 0.042929f
C13972 a_13623_n4162.t36 VSS 0.042774f
C13973 a_13623_n4162.t28 VSS 0.042774f
C13974 a_13623_n4162.t19 VSS 0.042774f
C13975 a_13623_n4162.t31 VSS 0.042774f
C13976 a_13623_n4162.t25 VSS 0.042774f
C13977 a_13623_n4162.t43 VSS 0.042774f
C13978 a_13623_n4162.t34 VSS 0.042774f
C13979 a_13623_n4162.t26 VSS 0.042774f
C13980 a_13623_n4162.t39 VSS 0.042774f
C13981 a_13623_n4162.t30 VSS 0.042794f
C13982 a_13623_n4162.t27 VSS 0.042937f
C13983 a_13623_n4162.t11 VSS 0.01101f
C13984 a_13623_n4162.t10 VSS 0.015244f
C13985 a_13623_n4162.n11 VSS 0.026254f
C13986 a_13623_n4162.n12 VSS 2.15567f
C13987 a_13623_n4162.n13 VSS 0.026583f
C13988 a_13623_n4162.t15 VSS 0.015244f
C13989 a_21772_1116.n0 VSS 0.588053f
C13990 a_21772_1116.t1 VSS 0.052911f
C13991 a_21772_1116.t2 VSS 0.058323f
C13992 a_21772_1116.t0 VSS 0.07776f
C13993 a_21772_1116.t3 VSS 0.065058f
C13994 a_21772_1116.t5 VSS 0.058056f
C13995 a_21772_1116.t13 VSS 0.055202f
C13996 a_21772_1116.n1 VSS 0.090091f
C13997 a_21772_1116.t17 VSS 0.058056f
C13998 a_21772_1116.t8 VSS 0.055202f
C13999 a_21772_1116.n2 VSS 0.090091f
C14000 a_21772_1116.t16 VSS 0.058056f
C14001 a_21772_1116.t6 VSS 0.055202f
C14002 a_21772_1116.n3 VSS -0.035108f
C14003 a_21772_1116.t4 VSS 0.058056f
C14004 a_21772_1116.t12 VSS 0.055202f
C14005 a_21772_1116.n4 VSS 0.101689f
C14006 a_21772_1116.t18 VSS 0.058056f
C14007 a_21772_1116.t9 VSS 0.055202f
C14008 a_21772_1116.n5 VSS 0.101689f
C14009 a_21772_1116.t15 VSS 0.058056f
C14010 a_21772_1116.t7 VSS 0.055202f
C14011 a_21772_1116.n6 VSS 0.101689f
C14012 a_21772_1116.t14 VSS 0.058056f
C14013 a_21772_1116.t11 VSS 0.055202f
C14014 a_21772_1116.n7 VSS 0.101689f
C14015 a_21772_1116.t19 VSS 0.058056f
C14016 a_21772_1116.t10 VSS 0.055202f
C14017 a_2167_3472.n0 VSS 3.15061f
C14018 a_2167_3472.t44 VSS 1.17475f
C14019 a_2167_3472.t58 VSS 1.09212f
C14020 a_2167_3472.t59 VSS 1.17326f
C14021 a_2167_3472.t27 VSS 1.0951f
C14022 a_2167_3472.t12 VSS 1.17178f
C14023 a_2167_3472.t70 VSS 1.09361f
C14024 a_2167_3472.t47 VSS 1.17326f
C14025 a_2167_3472.t79 VSS 1.17326f
C14026 a_2167_3472.t30 VSS 1.17178f
C14027 a_2167_3472.t25 VSS 1.17326f
C14028 a_2167_3472.t49 VSS 1.17178f
C14029 a_2167_3472.t65 VSS 1.17475f
C14030 a_2167_3472.t64 VSS 1.17178f
C14031 a_2167_3472.t11 VSS 1.17326f
C14032 a_2167_3472.t53 VSS 1.17178f
C14033 a_2167_3472.t57 VSS 1.09212f
C14034 a_2167_3472.t29 VSS 1.17178f
C14035 a_2167_3472.t23 VSS 1.17178f
C14036 a_2167_3472.t15 VSS 1.17178f
C14037 a_2167_3472.t76 VSS 1.17326f
C14038 a_2167_3472.t13 VSS 1.17178f
C14039 a_2167_3472.t20 VSS 1.01247f
C14040 a_2167_3472.t21 VSS 1.09361f
C14041 a_2167_3472.t22 VSS 1.09659f
C14042 a_2167_3472.t41 VSS 1.17475f
C14043 a_2167_3472.t73 VSS 1.09212f
C14044 a_2167_3472.t62 VSS 1.0951f
C14045 a_2167_3472.t50 VSS 1.0951f
C14046 a_2167_3472.t51 VSS 1.09212f
C14047 a_2167_3472.t66 VSS 1.09212f
C14048 a_2167_3472.t42 VSS 1.09361f
C14049 a_2167_3472.t45 VSS 1.01395f
C14050 a_2167_3472.t54 VSS 1.0951f
C14051 a_2167_3472.t71 VSS 1.17326f
C14052 a_2167_3472.t75 VSS 1.17624f
C14053 a_2167_3472.t14 VSS 1.17624f
C14054 a_2167_3472.t43 VSS 1.17326f
C14055 a_2167_3472.t83 VSS 1.17178f
C14056 a_2167_3472.t82 VSS 1.17326f
C14057 a_2167_3472.t60 VSS 1.17326f
C14058 a_2167_3472.t10 VSS 1.17326f
C14059 a_2167_3472.t77 VSS 1.17326f
C14060 a_2167_3472.t28 VSS 1.09659f
C14061 a_2167_3472.t52 VSS 1.09212f
C14062 a_2167_3472.t24 VSS 1.09361f
C14063 a_2167_3472.t18 VSS 1.09361f
C14064 a_2167_3472.t63 VSS 1.09212f
C14065 a_2167_3472.t67 VSS 1.01395f
C14066 a_2167_3472.t55 VSS 1.09361f
C14067 a_2167_3472.t69 VSS 1.09361f
C14068 a_2167_3472.t56 VSS 1.09361f
C14069 a_2167_3472.t46 VSS 1.09212f
C14070 a_2167_3472.t61 VSS 1.09361f
C14071 a_2167_3472.t84 VSS 0.150933f
C14072 a_2167_3472.t39 VSS 0.135774f
C14073 a_2167_3472.t8 VSS 0.131857f
C14074 a_2167_3472.t3 VSS 0.017055f
C14075 a_2167_3472.t6 VSS 0.017055f
C14076 a_2167_3472.n1 VSS 0.093873f
C14077 a_2167_3472.t34 VSS 0.017055f
C14078 a_2167_3472.t37 VSS 0.017055f
C14079 a_2167_3472.n2 VSS 0.091618f
C14080 a_2167_3472.t9 VSS 0.017055f
C14081 a_2167_3472.t2 VSS 0.017055f
C14082 a_2167_3472.n3 VSS 0.093558f
C14083 a_2167_3472.t40 VSS 0.017055f
C14084 a_2167_3472.t33 VSS 0.017055f
C14085 a_2167_3472.n4 VSS 0.092207f
C14086 a_2167_3472.t36 VSS 0.017055f
C14087 a_2167_3472.t31 VSS 0.017055f
C14088 a_2167_3472.n5 VSS 0.092207f
C14089 a_2167_3472.t5 VSS 0.017055f
C14090 a_2167_3472.t0 VSS 0.017055f
C14091 a_2167_3472.n6 VSS 0.093323f
C14092 a_2167_3472.t4 VSS 0.017055f
C14093 a_2167_3472.t7 VSS 0.017055f
C14094 a_2167_3472.n7 VSS 0.093401f
C14095 a_2167_3472.t35 VSS 0.017055f
C14096 a_2167_3472.t38 VSS 0.017055f
C14097 a_2167_3472.n8 VSS 0.091683f
C14098 a_2167_3472.t1 VSS 0.133274f
C14099 a_2167_3472.t32 VSS 0.135654f
C14100 a_2167_3472.n9 VSS 7.6709f
C14101 a_2167_3472.t19 VSS 1.15027f
C14102 a_2167_3472.t74 VSS 1.0951f
C14103 a_2167_3472.t68 VSS 1.17326f
C14104 a_2167_3472.t48 VSS 1.17326f
C14105 a_2167_3472.t78 VSS 1.17475f
C14106 a_2167_3472.t81 VSS 1.17475f
C14107 a_2167_3472.t26 VSS 1.17475f
C14108 a_2167_3472.t17 VSS 1.17475f
C14109 a_2167_3472.t16 VSS 1.17475f
C14110 a_2167_3472.t80 VSS 1.17178f
C14111 a_2167_3472.t72 VSS 1.17178f
C14112 a_11087_n23528.t39 VSS 0.933815f
C14113 a_11087_n23528.n0 VSS 1.20465f
C14114 a_11087_n23528.t60 VSS 0.933815f
C14115 a_11087_n23528.n1 VSS 1.33628f
C14116 a_11087_n23528.t44 VSS 2.44091f
C14117 a_11087_n23528.t35 VSS 2.18635f
C14118 a_11087_n23528.t57 VSS 0.933815f
C14119 a_11087_n23528.n2 VSS 1.35628f
C14120 a_11087_n23528.t49 VSS 0.933815f
C14121 a_11087_n23528.n3 VSS 0.691757f
C14122 a_11087_n23528.n4 VSS 0.403775f
C14123 a_11087_n23528.t38 VSS 1.88066f
C14124 a_11087_n23528.n5 VSS 0.050836f
C14125 a_11087_n23528.t50 VSS 1.94149f
C14126 a_11087_n23528.n6 VSS 0.248726f
C14127 a_11087_n23528.t53 VSS 1.98706f
C14128 a_11087_n23528.n7 VSS 0.360929f
C14129 a_11087_n23528.t52 VSS 0.933815f
C14130 a_11087_n23528.n8 VSS 0.933929f
C14131 a_11087_n23528.n9 VSS 0.365198f
C14132 a_11087_n23528.t48 VSS 0.933815f
C14133 a_11087_n23528.n10 VSS 0.813944f
C14134 a_11087_n23528.t56 VSS 0.933815f
C14135 a_11087_n23528.n11 VSS 0.813916f
C14136 a_11087_n23528.n12 VSS 0.466664f
C14137 a_11087_n23528.t47 VSS 0.933815f
C14138 a_11087_n23528.n13 VSS 0.818343f
C14139 a_11087_n23528.n14 VSS 0.360929f
C14140 a_11087_n23528.t30 VSS 0.933815f
C14141 a_11087_n23528.n15 VSS 0.857281f
C14142 a_11087_n23528.t32 VSS 0.933815f
C14143 a_11087_n23528.n16 VSS 0.05096f
C14144 a_11087_n23528.n17 VSS 0.925748f
C14145 a_11087_n23528.t45 VSS 0.933815f
C14146 a_11087_n23528.n18 VSS 0.117698f
C14147 a_11087_n23528.n19 VSS 0.050836f
C14148 a_11087_n23528.n20 VSS 0.8921f
C14149 a_11087_n23528.n21 VSS 0.033933f
C14150 a_11087_n23528.n22 VSS 0.032644f
C14151 a_11087_n23528.n23 VSS 0.095093f
C14152 a_11087_n23528.n24 VSS 0.033087f
C14153 a_11087_n23528.n25 VSS 0.032852f
C14154 a_11087_n23528.n26 VSS 0.03296f
C14155 a_11087_n23528.n27 VSS 0.032876f
C14156 a_11087_n23528.n28 VSS 0.033087f
C14157 a_11087_n23528.n29 VSS 0.089332f
C14158 a_11087_n23528.n30 VSS 0.033403f
C14159 a_11087_n23528.n31 VSS 0.032433f
C14160 a_11087_n23528.n32 VSS 0.112277f
C14161 a_11087_n23528.n33 VSS 0.032247f
C14162 a_11087_n23528.n34 VSS 0.038371f
C14163 a_11087_n23528.n35 VSS 0.0326f
C14164 a_11087_n23528.n36 VSS 0.038728f
C14165 a_11087_n23528.n37 VSS 0.032247f
C14166 a_11087_n23528.n38 VSS 0.067621f
C14167 a_11087_n23528.n39 VSS 0.139053f
C14168 a_11087_n23528.t55 VSS 1.77901f
C14169 a_11087_n23528.t37 VSS 1.73804f
C14170 a_11087_n23528.t41 VSS 1.74543f
C14171 a_11087_n23528.t46 VSS 1.9356f
C14172 a_11087_n23528.t33 VSS 1.95503f
C14173 a_11087_n23528.t43 VSS 1.73498f
C14174 a_11087_n23528.t61 VSS 1.65694f
C14175 a_11087_n23528.t58 VSS 2.0135f
C14176 a_11087_n23528.n52 VSS 0.167851f
C14177 a_11087_n23528.n56 VSS 0.123258f
C14178 a_11087_n23528.n58 VSS 0.013796f
C14179 a_11087_n23528.n59 VSS 0.013796f
C14180 a_11087_n23528.n64 VSS 0.03434f
C14181 a_11087_n23528.n65 VSS 0.03434f
C14182 a_11087_n23528.n70 VSS 0.013777f
C14183 a_11087_n23528.n71 VSS 0.013777f
C14184 a_11087_n23528.n76 VSS 0.034359f
C14185 a_11087_n23528.n77 VSS 0.034359f
C14186 a_11087_n23528.n82 VSS 0.013777f
C14187 a_11087_n23528.n83 VSS 0.013777f
C14188 a_11087_n23528.n88 VSS 0.031113f
C14189 a_11087_n23528.t31 VSS 1.9438f
C14190 a_11087_n23528.t59 VSS 1.73804f
C14191 a_11087_n23528.t40 VSS 1.80796f
C14192 a_11087_n23528.t51 VSS 1.95503f
C14193 a_11087_n23528.t36 VSS 1.9356f
C14194 a_11087_n23528.n101 VSS 0.071535f
C14195 a_11087_n23528.n106 VSS 0.013796f
C14196 a_11087_n23528.n107 VSS 0.013796f
C14197 a_11087_n23528.n112 VSS 0.034359f
C14198 a_11087_n23528.n113 VSS 0.034359f
C14199 a_11087_n23528.n118 VSS 0.013777f
C14200 a_11087_n23528.n119 VSS 0.013777f
C14201 a_11087_n23528.n124 VSS 0.091532f
C14202 a_11087_n23528.n125 VSS 0.091532f
C14203 a_11087_n23528.t42 VSS 1.62863f
C14204 a_11087_n23528.t34 VSS 1.80305f
C14205 a_11087_n23528.t54 VSS 2.04374f
C14206 a_11087_n23528.n130 VSS 0.013777f
C14207 a_11087_n23528.n131 VSS 0.013777f
C14208 a_11087_n23528.n136 VSS 0.675925f
C14209 a_11087_n23528.n137 VSS 0.780073f
C14210 a_11087_n23528.n138 VSS 0.033173f
C14211 a_11087_n23528.n139 VSS 0.15103f
C14212 a_11087_n23528.n140 VSS 0.033173f
C14213 a_11087_n23528.n141 VSS 0.033259f
C14214 a_11087_n23528.n142 VSS 0.032604f
C14215 a_11087_n23528.n143 VSS 0.032965f
C14216 a_11087_n23528.n144 VSS 0.032604f
C14217 a_11087_n23528.n145 VSS 0.033136f
C14218 a_11087_n23528.n146 VSS 0.044924f
C14219 a_11087_n23528.n147 VSS 0.032604f
C14220 a_22444_332.t19 VSS 0.862586f
C14221 a_22444_332.n0 VSS 1.21712f
C14222 a_22444_332.t26 VSS 0.444527f
C14223 a_22444_332.t15 VSS 0.109071f
C14224 a_22444_332.t1 VSS 2.41412f
C14225 a_22444_332.t3 VSS 0.087093f
C14226 a_22444_332.t5 VSS 0.094861f
C14227 a_22444_332.t4 VSS 0.102496f
C14228 a_22444_332.t6 VSS 0.030214f
C14229 a_22444_332.n1 VSS 1.26428f
C14230 a_22444_332.t0 VSS 0.045683f
C14231 a_22444_332.t2 VSS 0.107233f
C14232 a_22444_332.t8 VSS 0.054639f
C14233 a_22444_332.t21 VSS 0.062389f
C14234 a_22444_332.n2 VSS 0.08609f
C14235 a_22444_332.t22 VSS 0.062435f
C14236 a_22444_332.t12 VSS 0.064013f
C14237 a_22444_332.t32 VSS 0.055598f
C14238 a_22444_332.n3 VSS 0.075734f
C14239 a_22444_332.t11 VSS 0.068581f
C14240 a_22444_332.t14 VSS 0.051955f
C14241 a_22444_332.t20 VSS 0.063848f
C14242 a_22444_332.n4 VSS 0.452951f
C14243 a_22444_332.t34 VSS 0.026513f
C14244 a_22444_332.t33 VSS 0.02736f
C14245 a_22444_332.t36 VSS 0.062389f
C14246 a_22444_332.t7 VSS 0.054639f
C14247 a_22444_332.n5 VSS 0.115953f
C14248 a_22444_332.t31 VSS 0.028707f
C14249 a_22444_332.t27 VSS 0.191574f
C14250 a_22444_332.t13 VSS 0.052647f
C14251 a_22444_332.t29 VSS 0.06087f
C14252 a_22444_332.n6 VSS 0.265316f
C14253 a_22444_332.n7 VSS 0.584046f
C14254 a_22444_332.t25 VSS 0.02736f
C14255 a_22444_332.t18 VSS 0.02736f
C14256 a_22444_332.t10 VSS 0.115749f
C14257 a_22444_332.n8 VSS 0.948934f
C14258 a_22444_332.t24 VSS 0.026513f
C14259 a_22444_332.t16 VSS 0.120758f
C14260 a_22444_332.t17 VSS 0.052647f
C14261 a_22444_332.t23 VSS 0.06087f
C14262 a_22444_332.n9 VSS 0.113773f
C14263 a_22444_332.n10 VSS 0.581194f
C14264 a_22444_332.t35 VSS 0.02926f
C14265 a_22444_332.t9 VSS 0.026227f
C14266 a_22444_332.n11 VSS 0.1126f
C14267 a_22444_332.t28 VSS 0.052647f
C14268 a_22444_332.t30 VSS 0.06087f
C14269 a_22444_332.n12 VSS 0.146859f
C14270 a_22444_332.n13 VSS 1.30092f
C14271 a_22444_332.n14 VSS 1.44792f
C14272 EOC.t11 VSS 0.034759f
C14273 EOC.t10 VSS 0.025104f
C14274 EOC.n0 VSS 0.060614f
C14275 EOC.t9 VSS 0.034759f
C14276 EOC.t15 VSS 0.025104f
C14277 EOC.n1 VSS 0.076677f
C14278 EOC.n2 VSS 0.189109f
C14279 EOC.t13 VSS 0.034759f
C14280 EOC.t12 VSS 0.025104f
C14281 EOC.n3 VSS 0.060614f
C14282 EOC.t8 VSS 0.025104f
C14283 EOC.t14 VSS 0.034759f
C14284 EOC.n4 VSS 0.075598f
C14285 EOC.n5 VSS 0.190187f
C14286 EOC.t1 VSS 0.016873f
C14287 EOC.t0 VSS 0.016873f
C14288 EOC.n6 VSS 0.033863f
C14289 EOC.t4 VSS 0.016873f
C14290 EOC.t2 VSS 0.016873f
C14291 EOC.n7 VSS 0.040715f
C14292 EOC.n8 VSS 0.182121f
C14293 EOC.t7 VSS 0.016873f
C14294 EOC.t6 VSS 0.016873f
C14295 EOC.n9 VSS 0.033863f
C14296 EOC.t5 VSS 0.016873f
C14297 EOC.t3 VSS 0.016873f
C14298 EOC.n10 VSS 0.04058f
C14299 EOC.n11 VSS 0.185334f
C14300 EOC.n12 VSS 0.149041f
C14301 EOC.n13 VSS 0.132801f
C14302 EOC.n14 VSS 0.232613f
C14303 a_45648_1564.n0 VSS 0.383346f
C14304 a_45648_1564.t5 VSS 0.019652f
C14305 a_45648_1564.t6 VSS 0.027211f
C14306 a_45648_1564.t4 VSS 0.019652f
C14307 a_45648_1564.n1 VSS 0.047321f
C14308 a_45648_1564.t3 VSS 0.013209f
C14309 a_45648_1564.t1 VSS 0.013209f
C14310 a_45648_1564.n2 VSS 0.026494f
C14311 a_45648_1564.t0 VSS 0.013209f
C14312 a_45648_1564.t2 VSS 0.013209f
C14313 a_45648_1564.n3 VSS 0.031906f
C14314 a_45648_1564.t17 VSS 0.058056f
C14315 a_45648_1564.t14 VSS 0.055202f
C14316 a_45648_1564.n4 VSS 0.090091f
C14317 a_45648_1564.t9 VSS 0.058056f
C14318 a_45648_1564.t19 VSS 0.055202f
C14319 a_45648_1564.n5 VSS -0.035108f
C14320 a_45648_1564.t15 VSS 0.058056f
C14321 a_45648_1564.t8 VSS 0.055202f
C14322 a_45648_1564.n6 VSS 0.101689f
C14323 a_45648_1564.t16 VSS 0.058056f
C14324 a_45648_1564.t11 VSS 0.055202f
C14325 a_45648_1564.n7 VSS 0.101689f
C14326 a_45648_1564.t12 VSS 0.058056f
C14327 a_45648_1564.t21 VSS 0.055202f
C14328 a_45648_1564.n8 VSS 0.101689f
C14329 a_45648_1564.t13 VSS 0.058056f
C14330 a_45648_1564.t23 VSS 0.055202f
C14331 a_45648_1564.n9 VSS 0.101689f
C14332 a_45648_1564.t10 VSS 0.058056f
C14333 a_45648_1564.t20 VSS 0.055202f
C14334 a_45648_1564.n10 VSS 0.090091f
C14335 a_45648_1564.t22 VSS 0.058056f
C14336 a_45648_1564.t18 VSS 0.055202f
C14337 a_45648_1564.n11 VSS 0.146257f
C14338 a_45648_1564.n12 VSS 0.060222f
C14339 a_45648_1564.t7 VSS 0.027211f
C14340 a_24815_n3588.n0 VSS 0.920329f
C14341 a_24815_n3588.t0 VSS 0.074613f
C14342 a_24815_n3588.n1 VSS 0.181232f
C14343 a_24815_n3588.n3 VSS 0.181232f
C14344 a_24815_n3588.n4 VSS 0.576962f
C14345 a_24815_n3588.t3 VSS 0.964165f
C14346 a_24815_n3588.t2 VSS 0.15329f
C14347 a_24815_n3588.t1 VSS 0.041326f
C14348 a_24815_n3588.t11 VSS 0.07614f
C14349 a_24815_n3588.t22 VSS 0.069899f
C14350 a_24815_n3588.n5 VSS 0.210668f
C14351 a_24815_n3588.t18 VSS 0.132457f
C14352 a_24815_n3588.t23 VSS 0.089828f
C14353 a_24815_n3588.n6 VSS 0.151063f
C14354 a_24815_n3588.t13 VSS 0.107561f
C14355 a_24815_n3588.t4 VSS 0.118805f
C14356 a_24815_n3588.n7 VSS 0.157301f
C14357 a_24815_n3588.t10 VSS 0.087573f
C14358 a_24815_n3588.t17 VSS 0.116817f
C14359 a_24815_n3588.n8 VSS 0.240001f
C14360 a_24815_n3588.t6 VSS 0.10108f
C14361 a_24815_n3588.t5 VSS 0.116179f
C14362 a_24815_n3588.n9 VSS 0.394824f
C14363 a_24815_n3588.t12 VSS 0.116498f
C14364 a_24815_n3588.t21 VSS 0.10108f
C14365 a_24815_n3588.n10 VSS 0.49827f
C14366 a_24815_n3588.n11 VSS 2.19353f
C14367 a_24815_n3588.n12 VSS 1.51907f
C14368 a_24815_n3588.t7 VSS 0.098305f
C14369 a_24815_n3588.t14 VSS 0.127539f
C14370 a_24815_n3588.n13 VSS 0.188757f
C14371 a_24815_n3588.t15 VSS 0.098305f
C14372 a_24815_n3588.t20 VSS 0.098305f
C14373 a_24815_n3588.t16 VSS 0.115676f
C14374 a_24815_n3588.t19 VSS 0.115676f
C14375 a_24815_n3588.t9 VSS 0.098305f
C14376 a_24815_n3588.t8 VSS 0.127597f
C14377 a_24815_n3588.n14 VSS 0.154042f
C14378 a_24815_n3588.n15 VSS 0.800368f
C14379 a_24815_n3588.n16 VSS 1.28533f
C14380 a_21692_n6694.t1 VSS 0.126336f
C14381 a_21692_n6694.t0 VSS 0.077364f
C14382 a_21692_n6694.n0 VSS 0.699732f
C14383 a_21692_n6694.n1 VSS 1.31156f
C14384 a_21692_n6694.t16 VSS 0.033832f
C14385 a_21692_n6694.t12 VSS 0.03702f
C14386 a_21692_n6694.n2 VSS 0.290796f
C14387 a_21692_n6694.t20 VSS 0.050579f
C14388 a_21692_n6694.t34 VSS 0.084884f
C14389 a_21692_n6694.n3 VSS 0.146713f
C14390 a_21692_n6694.n4 VSS 0.833285f
C14391 a_21692_n6694.t6 VSS 0.037734f
C14392 a_21692_n6694.t8 VSS 0.033822f
C14393 a_21692_n6694.n5 VSS 0.094152f
C14394 a_21692_n6694.t19 VSS 0.075406f
C14395 a_21692_n6694.t15 VSS 0.056293f
C14396 a_21692_n6694.n6 VSS 0.320777f
C14397 a_21692_n6694.t9 VSS 0.079447f
C14398 a_21692_n6694.t14 VSS 0.072934f
C14399 a_21692_n6694.n7 VSS 0.145069f
C14400 a_21692_n6694.n8 VSS 1.39765f
C14401 a_21692_n6694.n9 VSS 0.420022f
C14402 a_21692_n6694.t13 VSS 0.037734f
C14403 a_21692_n6694.t17 VSS 0.033822f
C14404 a_21692_n6694.n10 VSS 0.094152f
C14405 a_21692_n6694.n11 VSS 0.480628f
C14406 a_21692_n6694.t5 VSS 0.08073f
C14407 a_21692_n6694.t31 VSS 0.069305f
C14408 a_21692_n6694.n12 VSS 0.096498f
C14409 a_21692_n6694.t27 VSS 0.082537f
C14410 a_21692_n6694.t35 VSS 0.063869f
C14411 a_21692_n6694.n13 VSS 0.094647f
C14412 a_21692_n6694.n14 VSS 0.283834f
C14413 a_21692_n6694.n15 VSS 0.273526f
C14414 a_21692_n6694.t11 VSS 0.033832f
C14415 a_21692_n6694.t10 VSS 0.03702f
C14416 a_21692_n6694.n16 VSS 0.121462f
C14417 a_21692_n6694.t32 VSS 0.03702f
C14418 a_21692_n6694.t25 VSS 0.033832f
C14419 a_21692_n6694.n17 VSS 0.124232f
C14420 a_21692_n6694.t3 VSS 0.067893f
C14421 a_21692_n6694.t7 VSS 0.078497f
C14422 a_21692_n6694.n18 VSS 0.164034f
C14423 a_21692_n6694.t21 VSS 0.033832f
C14424 a_21692_n6694.t18 VSS 0.03702f
C14425 a_21692_n6694.n19 VSS 0.17508f
C14426 a_21692_n6694.t26 VSS 0.03702f
C14427 a_21692_n6694.t23 VSS 0.033832f
C14428 a_21692_n6694.n20 VSS 0.101701f
C14429 a_21692_n6694.n21 VSS 0.282246f
C14430 a_21692_n6694.t24 VSS 0.079447f
C14431 a_21692_n6694.t33 VSS 0.072934f
C14432 a_21692_n6694.n22 VSS 0.100151f
C14433 a_21692_n6694.n23 VSS 0.478402f
C14434 a_21692_n6694.t29 VSS 0.037734f
C14435 a_21692_n6694.t28 VSS 0.033822f
C14436 a_21692_n6694.n24 VSS 0.696547f
C14437 a_21692_n6694.t2 VSS 0.065248f
C14438 a_21692_n6694.t4 VSS 0.074994f
C14439 a_21692_n6694.n25 VSS 0.118371f
C14440 a_21692_n6694.n26 VSS 0.499383f
C14441 a_21692_n6694.t22 VSS 0.064652f
C14442 a_21692_n6694.t30 VSS 0.06016f
C14443 a_21692_n6694.n27 VSS 0.151394f
C14444 a_21692_n6694.n28 VSS 0.776253f
C14445 a_21692_n6694.n29 VSS 0.589742f
C14446 a_21692_n6694.n30 VSS 0.666919f
C14447 a_21692_n6694.n31 VSS 0.218605f
C14448 a_13623_n6840.n0 VSS 3.65914f
C14449 a_13623_n6840.n1 VSS 5.54012f
C14450 a_13623_n6840.n2 VSS 0.474608f
C14451 a_13623_n6840.n3 VSS 0.084524f
C14452 a_13623_n6840.n4 VSS 0.319233f
C14453 a_13623_n6840.t9 VSS 0.011651f
C14454 a_13623_n6840.t12 VSS 0.011651f
C14455 a_13623_n6840.t13 VSS 0.016132f
C14456 a_13623_n6840.n5 VSS 0.028131f
C14457 a_13623_n6840.t10 VSS 0.011651f
C14458 a_13623_n6840.t14 VSS 0.016132f
C14459 a_13623_n6840.n6 VSS 0.028131f
C14460 a_13623_n6840.t8 VSS 0.011651f
C14461 a_13623_n6840.t11 VSS 0.016132f
C14462 a_13623_n6840.n7 VSS 0.028131f
C14463 a_13623_n6840.t38 VSS 0.045265f
C14464 a_13623_n6840.t20 VSS 0.045438f
C14465 a_13623_n6840.t26 VSS 0.045265f
C14466 a_13623_n6840.t36 VSS 0.045438f
C14467 a_13623_n6840.t31 VSS 0.045265f
C14468 a_13623_n6840.t41 VSS 0.045438f
C14469 a_13623_n6840.t16 VSS 0.045265f
C14470 a_13623_n6840.t23 VSS 0.045265f
C14471 a_13623_n6840.t33 VSS 0.045265f
C14472 a_13623_n6840.t19 VSS 0.045265f
C14473 a_13623_n6840.t27 VSS 0.045265f
C14474 a_13623_n6840.t40 VSS 0.045265f
C14475 a_13623_n6840.t30 VSS 0.045523f
C14476 a_13623_n6840.t39 VSS 0.04543f
C14477 a_13623_n6840.t22 VSS 0.045265f
C14478 a_13623_n6840.t45 VSS 0.045265f
C14479 a_13623_n6840.t35 VSS 0.045265f
C14480 a_13623_n6840.t18 VSS 0.045265f
C14481 a_13623_n6840.t42 VSS 0.045265f
C14482 a_13623_n6840.t28 VSS 0.045265f
C14483 a_13623_n6840.t21 VSS 0.045265f
C14484 a_13623_n6840.t43 VSS 0.045265f
C14485 a_13623_n6840.t24 VSS 0.045265f
C14486 a_13623_n6840.t17 VSS 0.045287f
C14487 a_13623_n6840.t25 VSS 0.045438f
C14488 a_13623_n6840.t37 VSS 0.045438f
C14489 a_13623_n6840.t32 VSS 0.045438f
C14490 a_13623_n6840.t44 VSS 0.045438f
C14491 a_13623_n6840.t34 VSS 0.045438f
C14492 a_13623_n6840.t29 VSS 0.045438f
C14493 a_13623_n6840.n8 VSS 0.015716f
C14494 a_13623_n6840.n9 VSS 0.018834f
C14495 a_13623_n6840.n10 VSS 0.015716f
C14496 a_13623_n6840.n11 VSS 0.018896f
C14497 a_13623_n6840.n12 VSS 0.035086f
C14498 a_13623_n6840.t15 VSS 0.016132f
C14499 a_21772_n20836.n0 VSS 0.400111f
C14500 a_21772_n20836.t4 VSS 0.020507f
C14501 a_21772_n20836.t6 VSS 0.020507f
C14502 a_21772_n20836.t5 VSS 0.028394f
C14503 a_21772_n20836.n1 VSS 0.049378f
C14504 a_21772_n20836.t3 VSS 0.013783f
C14505 a_21772_n20836.t2 VSS 0.013783f
C14506 a_21772_n20836.n2 VSS 0.027645f
C14507 a_21772_n20836.t1 VSS 0.013783f
C14508 a_21772_n20836.t0 VSS 0.013783f
C14509 a_21772_n20836.n3 VSS 0.033293f
C14510 a_21772_n20836.t8 VSS 0.06058f
C14511 a_21772_n20836.t16 VSS 0.057602f
C14512 a_21772_n20836.n4 VSS 0.094008f
C14513 a_21772_n20836.t20 VSS 0.06058f
C14514 a_21772_n20836.t13 VSS 0.057602f
C14515 a_21772_n20836.n5 VSS 0.094008f
C14516 a_21772_n20836.t23 VSS 0.06058f
C14517 a_21772_n20836.t10 VSS 0.057602f
C14518 a_21772_n20836.n6 VSS -0.036634f
C14519 a_21772_n20836.t9 VSS 0.06058f
C14520 a_21772_n20836.t17 VSS 0.057602f
C14521 a_21772_n20836.n7 VSS 0.106111f
C14522 a_21772_n20836.t21 VSS 0.06058f
C14523 a_21772_n20836.t14 VSS 0.057602f
C14524 a_21772_n20836.n8 VSS 0.106111f
C14525 a_21772_n20836.t18 VSS 0.06058f
C14526 a_21772_n20836.t11 VSS 0.057602f
C14527 a_21772_n20836.n9 VSS 0.106111f
C14528 a_21772_n20836.t19 VSS 0.06058f
C14529 a_21772_n20836.t12 VSS 0.057602f
C14530 a_21772_n20836.n10 VSS 0.106111f
C14531 a_21772_n20836.t22 VSS 0.06058f
C14532 a_21772_n20836.t15 VSS 0.057602f
C14533 a_21772_n20836.n11 VSS 0.152518f
C14534 a_21772_n20836.n12 VSS 0.06284f
C14535 a_21772_n20836.t7 VSS 0.028394f
C14536 a_11087_n12816.t3 VSS 0.026453f
C14537 a_11087_n12816.t15 VSS 0.026453f
C14538 a_11087_n12816.t13 VSS 0.026453f
C14539 a_11087_n12816.n0 VSS 0.129398f
C14540 a_11087_n12816.t17 VSS 0.026453f
C14541 a_11087_n12816.t10 VSS 0.026453f
C14542 a_11087_n12816.n1 VSS 0.124481f
C14543 a_11087_n12816.n2 VSS 0.362621f
C14544 a_11087_n12816.t14 VSS 0.026453f
C14545 a_11087_n12816.t18 VSS 0.026453f
C14546 a_11087_n12816.n3 VSS 0.126171f
C14547 a_11087_n12816.n4 VSS 0.125275f
C14548 a_11087_n12816.t11 VSS 0.026453f
C14549 a_11087_n12816.t19 VSS 0.026453f
C14550 a_11087_n12816.n5 VSS 0.125688f
C14551 a_11087_n12816.n6 VSS 0.125369f
C14552 a_11087_n12816.t12 VSS 0.026453f
C14553 a_11087_n12816.t16 VSS 0.026453f
C14554 a_11087_n12816.n7 VSS 0.126171f
C14555 a_11087_n12816.n8 VSS 0.340653f
C14556 a_11087_n12816.t23 VSS 0.026453f
C14557 a_11087_n12816.t25 VSS 0.026453f
C14558 a_11087_n12816.n9 VSS 0.127376f
C14559 a_11087_n12816.t21 VSS 0.026453f
C14560 a_11087_n12816.t28 VSS 0.026453f
C14561 a_11087_n12816.n10 VSS 0.123678f
C14562 a_11087_n12816.n11 VSS 0.42815f
C14563 a_11087_n12816.t24 VSS 0.026453f
C14564 a_11087_n12816.t20 VSS 0.026453f
C14565 a_11087_n12816.n12 VSS 0.122969f
C14566 a_11087_n12816.n13 VSS 0.146322f
C14567 a_11087_n12816.t27 VSS 0.026453f
C14568 a_11087_n12816.t29 VSS 0.026453f
C14569 a_11087_n12816.n14 VSS 0.124315f
C14570 a_11087_n12816.n15 VSS 0.147681f
C14571 a_11087_n12816.t26 VSS 0.026453f
C14572 a_11087_n12816.t22 VSS 0.026453f
C14573 a_11087_n12816.n16 VSS 0.122969f
C14574 a_11087_n12816.n17 VSS 0.257862f
C14575 a_11087_n12816.n18 VSS 0.530252f
C14576 a_11087_n12816.t4 VSS 0.026453f
C14577 a_11087_n12816.t7 VSS 0.026453f
C14578 a_11087_n12816.n19 VSS 0.12433f
C14579 a_11087_n12816.n20 VSS 0.171311f
C14580 a_11087_n12816.t1 VSS 0.026453f
C14581 a_11087_n12816.t8 VSS 0.026453f
C14582 a_11087_n12816.n21 VSS 0.12433f
C14583 a_11087_n12816.n22 VSS 0.12636f
C14584 a_11087_n12816.t2 VSS 0.026453f
C14585 a_11087_n12816.t5 VSS 0.026453f
C14586 a_11087_n12816.n23 VSS 0.12433f
C14587 a_11087_n12816.n24 VSS 0.125706f
C14588 a_11087_n12816.t30 VSS 6.22367f
C14589 a_11087_n12816.t6 VSS 0.026453f
C14590 a_11087_n12816.t0 VSS 0.026453f
C14591 a_11087_n12816.n25 VSS 0.126499f
C14592 a_11087_n12816.n26 VSS 1.48916f
C14593 a_11087_n12816.n27 VSS 0.126829f
C14594 a_11087_n12816.n28 VSS 0.126499f
C14595 a_11087_n12816.t9 VSS 0.026453f
C14596 a_11023_n12196.n0 VSS 0.904871f
C14597 a_11023_n12196.t29 VSS 0.065212f
C14598 a_11023_n12196.n1 VSS 0.782917f
C14599 a_11023_n12196.n2 VSS 1.64085f
C14600 a_11023_n12196.t15 VSS 0.219126f
C14601 a_11023_n12196.t18 VSS 0.234136f
C14602 a_11023_n12196.t10 VSS 0.0377f
C14603 a_11023_n12196.t31 VSS 0.064062f
C14604 a_11023_n12196.t25 VSS 0.064062f
C14605 a_11023_n12196.t39 VSS 0.064062f
C14606 a_11023_n12196.t30 VSS 0.064062f
C14607 a_11023_n12196.t36 VSS 0.064062f
C14608 a_11023_n12196.t34 VSS 0.064062f
C14609 a_11023_n12196.t38 VSS 0.06392f
C14610 a_11023_n12196.t27 VSS 0.063818f
C14611 a_11023_n12196.t33 VSS 0.063818f
C14612 a_11023_n12196.t20 VSS 0.063818f
C14613 a_11023_n12196.t28 VSS 0.063818f
C14614 a_11023_n12196.t35 VSS 0.063818f
C14615 a_11023_n12196.t22 VSS 0.063818f
C14616 a_11023_n12196.t37 VSS 0.063818f
C14617 a_11023_n12196.t24 VSS 0.063818f
C14618 a_11023_n12196.t32 VSS 0.063818f
C14619 a_11023_n12196.t26 VSS 0.064062f
C14620 a_11023_n12196.t21 VSS 0.064062f
C14621 a_11023_n12196.t23 VSS 0.064062f
C14622 a_11023_n12196.t8 VSS 0.216709f
C14623 a_11023_n12196.t1 VSS 0.0377f
C14624 a_11023_n12196.t2 VSS 0.216709f
C14625 a_11023_n12196.t17 VSS 0.0377f
C14626 a_11023_n12196.t6 VSS 0.216709f
C14627 a_11023_n12196.t12 VSS 0.0377f
C14628 a_11023_n12196.t0 VSS 0.216709f
C14629 a_11023_n12196.t13 VSS 0.0377f
C14630 a_11023_n12196.t16 VSS 0.236521f
C14631 a_11023_n12196.t7 VSS 0.0377f
C14632 a_11023_n12196.n3 VSS 0.696191f
C14633 a_11023_n12196.n4 VSS 0.29804f
C14634 a_11023_n12196.n5 VSS 0.29804f
C14635 a_11023_n12196.n6 VSS 0.414463f
C14636 a_11023_n12196.n7 VSS 0.801546f
C14637 a_11023_n12196.t11 VSS 0.219124f
C14638 a_11023_n12196.t4 VSS 0.0377f
C14639 a_11023_n12196.n8 VSS 0.319464f
C14640 a_11023_n12196.t5 VSS 0.219124f
C14641 a_11023_n12196.t19 VSS 0.0377f
C14642 a_11023_n12196.n9 VSS 0.184638f
C14643 a_11023_n12196.t9 VSS 0.219124f
C14644 a_11023_n12196.t14 VSS 0.0377f
C14645 a_11023_n12196.n10 VSS 0.184638f
C14646 a_11023_n12196.n11 VSS 0.503296f
C14647 a_11023_n12196.t3 VSS 0.0377f
C14648 a_28156_n6412.n0 VSS 0.721559f
C14649 a_28156_n6412.n1 VSS 0.308352f
C14650 a_28156_n6412.n2 VSS 0.215117f
C14651 a_28156_n6412.t12 VSS 0.044777f
C14652 a_28156_n6412.t14 VSS 0.044777f
C14653 a_28156_n6412.t11 VSS 0.044777f
C14654 a_28156_n6412.n3 VSS 0.111909f
C14655 a_28156_n6412.t9 VSS 0.044777f
C14656 a_28156_n6412.t13 VSS 0.044777f
C14657 a_28156_n6412.n4 VSS 0.090675f
C14658 a_28156_n6412.t10 VSS 0.044777f
C14659 a_28156_n6412.t8 VSS 0.044777f
C14660 a_28156_n6412.n5 VSS 0.091938f
C14661 a_28156_n6412.t25 VSS 0.048019f
C14662 a_28156_n6412.t18 VSS 0.085014f
C14663 a_28156_n6412.n6 VSS 0.14664f
C14664 a_28156_n6412.t26 VSS 0.048019f
C14665 a_28156_n6412.t27 VSS 0.085014f
C14666 a_28156_n6412.n7 VSS 0.15398f
C14667 a_28156_n6412.t21 VSS 0.128938f
C14668 a_28156_n6412.t20 VSS 0.048019f
C14669 a_28156_n6412.t17 VSS 0.085014f
C14670 a_28156_n6412.n8 VSS 0.22715f
C14671 a_28156_n6412.n9 VSS 0.24834f
C14672 a_28156_n6412.t24 VSS 0.085014f
C14673 a_28156_n6412.t16 VSS 0.047713f
C14674 a_28156_n6412.n10 VSS 0.146945f
C14675 a_28156_n6412.t28 VSS 0.085014f
C14676 a_28156_n6412.t29 VSS 0.047713f
C14677 a_28156_n6412.n11 VSS 0.154286f
C14678 a_28156_n6412.t23 VSS 0.128938f
C14679 a_28156_n6412.t19 VSS 0.085014f
C14680 a_28156_n6412.t22 VSS 0.047713f
C14681 a_28156_n6412.n12 VSS 0.227455f
C14682 a_28156_n6412.n13 VSS 0.276729f
C14683 a_28156_n6412.n14 VSS 0.57208f
C14684 a_28156_n6412.t5 VSS 0.011398f
C14685 a_28156_n6412.t4 VSS 0.011398f
C14686 a_28156_n6412.n15 VSS 0.02315f
C14687 a_28156_n6412.t6 VSS 0.011398f
C14688 a_28156_n6412.t7 VSS 0.011398f
C14689 a_28156_n6412.n16 VSS 0.032657f
C14690 a_28156_n6412.t2 VSS 0.011398f
C14691 a_28156_n6412.t3 VSS 0.011398f
C14692 a_28156_n6412.n17 VSS 0.02315f
C14693 a_28156_n6412.t0 VSS 0.011398f
C14694 a_28156_n6412.t1 VSS 0.011398f
C14695 a_28156_n6412.n18 VSS 0.032657f
C14696 a_28156_n6412.n19 VSS 0.090675f
C14697 a_28156_n6412.t15 VSS 0.044777f
C14698 a_29800_n5940.n0 VSS 0.448816f
C14699 a_29800_n5940.t5 VSS 0.023188f
C14700 a_29800_n5940.t3 VSS 0.023188f
C14701 a_29800_n5940.t4 VSS 0.023188f
C14702 a_29800_n5940.n1 VSS 0.046856f
C14703 a_29800_n5940.t2 VSS 0.020552f
C14704 a_29800_n5940.n2 VSS 0.024427f
C14705 a_29800_n5940.t22 VSS 0.044539f
C14706 a_29800_n5940.t9 VSS 0.073413f
C14707 a_29800_n5940.n3 VSS 0.106957f
C14708 a_29800_n5940.t21 VSS 0.044539f
C14709 a_29800_n5940.t14 VSS 0.073413f
C14710 a_29800_n5940.n4 VSS 0.109926f
C14711 a_29800_n5940.t7 VSS 0.044539f
C14712 a_29800_n5940.t19 VSS 0.073413f
C14713 a_29800_n5940.n5 VSS 0.106957f
C14714 a_29800_n5940.t12 VSS 0.044539f
C14715 a_29800_n5940.t17 VSS 0.073413f
C14716 a_29800_n5940.n6 VSS -0.028686f
C14717 a_29800_n5940.t15 VSS 0.044539f
C14718 a_29800_n5940.t10 VSS 0.073413f
C14719 a_29800_n5940.n7 VSS 0.121662f
C14720 a_29800_n5940.t13 VSS 0.044539f
C14721 a_29800_n5940.t18 VSS 0.073413f
C14722 a_29800_n5940.n8 VSS 0.121662f
C14723 a_29800_n5940.t16 VSS 0.044539f
C14724 a_29800_n5940.t11 VSS 0.073413f
C14725 a_29800_n5940.n9 VSS 0.121662f
C14726 a_29800_n5940.t20 VSS 0.044539f
C14727 a_29800_n5940.t8 VSS 0.073413f
C14728 a_29800_n5940.n10 VSS 0.118692f
C14729 a_29800_n5940.n11 VSS 0.071373f
C14730 a_29800_n5940.n12 VSS 0.056236f
C14731 a_29800_n5940.t6 VSS 0.023188f
C14732 a_27884_332.t1 VSS 0.25015f
C14733 a_27884_332.t5 VSS 0.026344f
C14734 a_27884_332.t3 VSS 0.033868f
C14735 a_27884_332.n0 VSS 0.413971f
C14736 a_27884_332.t4 VSS 0.022363f
C14737 a_27884_332.t2 VSS 0.038469f
C14738 a_27884_332.n1 VSS 0.088933f
C14739 a_27884_332.n2 VSS 1.20414f
C14740 a_27884_332.t0 VSS 0.021759f
C14741 a_31628_n5940.n0 VSS 0.194444f
C14742 a_31628_n5940.n1 VSS 0.884727f
C14743 a_31628_n5940.n2 VSS 0.145504f
C14744 a_31628_n5940.t30 VSS 0.039743f
C14745 a_31628_n5940.t17 VSS 0.055029f
C14746 a_31628_n5940.t19 VSS 0.039743f
C14747 a_31628_n5940.n3 VSS 0.111732f
C14748 a_31628_n5940.t18 VSS 0.039743f
C14749 a_31628_n5940.t20 VSS 0.055029f
C14750 a_31628_n5940.n4 VSS 0.094772f
C14751 a_31628_n5940.n5 VSS 0.428611f
C14752 a_31628_n5940.t27 VSS 0.039743f
C14753 a_31628_n5940.t25 VSS 0.055029f
C14754 a_31628_n5940.n6 VSS 0.094772f
C14755 a_31628_n5940.n7 VSS 0.303087f
C14756 a_31628_n5940.t28 VSS 0.039743f
C14757 a_31628_n5940.t26 VSS 0.055029f
C14758 a_31628_n5940.n8 VSS 0.094772f
C14759 a_31628_n5940.t2 VSS 0.0158f
C14760 a_31628_n5940.t3 VSS 0.0158f
C14761 a_31628_n5940.n9 VSS 0.032025f
C14762 a_31628_n5940.t1 VSS 0.0158f
C14763 a_31628_n5940.t9 VSS 0.0158f
C14764 a_31628_n5940.n10 VSS 0.032025f
C14765 a_31628_n5940.t7 VSS 0.0158f
C14766 a_31628_n5940.t8 VSS 0.0158f
C14767 a_31628_n5940.n11 VSS 0.032025f
C14768 a_31628_n5940.t10 VSS 0.0158f
C14769 a_31628_n5940.t15 VSS 0.0158f
C14770 a_31628_n5940.n12 VSS 0.043516f
C14771 a_31628_n5940.n13 VSS 0.326828f
C14772 a_31628_n5940.n14 VSS 0.209454f
C14773 a_31628_n5940.t14 VSS 0.0158f
C14774 a_31628_n5940.t0 VSS 0.0158f
C14775 a_31628_n5940.n15 VSS 0.032025f
C14776 a_31628_n5940.t13 VSS 0.0158f
C14777 a_31628_n5940.t11 VSS 0.0158f
C14778 a_31628_n5940.n16 VSS 0.032025f
C14779 a_31628_n5940.t5 VSS 0.0158f
C14780 a_31628_n5940.t12 VSS 0.0158f
C14781 a_31628_n5940.n17 VSS 0.032025f
C14782 a_31628_n5940.t4 VSS 0.0158f
C14783 a_31628_n5940.t6 VSS 0.0158f
C14784 a_31628_n5940.n18 VSS 0.043516f
C14785 a_31628_n5940.n19 VSS 0.326828f
C14786 a_31628_n5940.n20 VSS 0.209454f
C14787 a_31628_n5940.t24 VSS 0.039743f
C14788 a_31628_n5940.t23 VSS 0.055029f
C14789 a_31628_n5940.n21 VSS 0.094828f
C14790 a_31628_n5940.t38 VSS 0.059014f
C14791 a_31628_n5940.t32 VSS 0.104479f
C14792 a_31628_n5940.n22 VSS 0.180215f
C14793 a_31628_n5940.t34 VSS 0.059014f
C14794 a_31628_n5940.t35 VSS 0.104479f
C14795 a_31628_n5940.n23 VSS 0.189236f
C14796 a_31628_n5940.t36 VSS 0.15846f
C14797 a_31628_n5940.t33 VSS 0.059014f
C14798 a_31628_n5940.t42 VSS 0.104479f
C14799 a_31628_n5940.n24 VSS 0.279159f
C14800 a_31628_n5940.n25 VSS 0.536317f
C14801 a_31628_n5940.t39 VSS 0.15846f
C14802 a_31628_n5940.t44 VSS 0.059014f
C14803 a_31628_n5940.t45 VSS 0.104479f
C14804 a_31628_n5940.n26 VSS 0.279159f
C14805 a_31628_n5940.t40 VSS 0.059014f
C14806 a_31628_n5940.t41 VSS 0.104479f
C14807 a_31628_n5940.n27 VSS 0.180215f
C14808 a_31628_n5940.t43 VSS 0.059014f
C14809 a_31628_n5940.t37 VSS 0.104479f
C14810 a_31628_n5940.n28 VSS 0.189236f
C14811 a_31628_n5940.n29 VSS 0.30297f
C14812 a_31628_n5940.n30 VSS 0.685657f
C14813 a_31628_n5940.n31 VSS 0.191129f
C14814 a_31628_n5940.t21 VSS 0.039743f
C14815 a_31628_n5940.t22 VSS 0.055029f
C14816 a_31628_n5940.n32 VSS 0.094772f
C14817 a_31628_n5940.n33 VSS 0.291459f
C14818 a_31628_n5940.t29 VSS 0.039743f
C14819 a_31628_n5940.t16 VSS 0.055029f
C14820 a_31628_n5940.n34 VSS 0.094772f
C14821 a_31628_n5940.n35 VSS 0.303087f
C14822 a_31628_n5940.n36 VSS 0.094772f
C14823 a_31628_n5940.t31 VSS 0.055029f
C14824 a_33496_n6659.n0 VSS 3.38274f
C14825 a_33496_n6659.t2 VSS 0.147698f
C14826 a_33496_n6659.t0 VSS 0.058719f
C14827 a_33496_n6659.t7 VSS 0.058719f
C14828 a_33496_n6659.t4 VSS 0.147698f
C14829 a_33496_n6659.t3 VSS 0.147698f
C14830 a_33496_n6659.n1 VSS 0.303673f
C14831 a_33496_n6659.n2 VSS 0.303673f
C14832 a_33496_n6659.t5 VSS 0.168139f
C14833 a_33496_n6659.t6 VSS 0.050967f
C14834 a_33496_n6659.t1 VSS 0.064596f
C14835 a_33496_n6659.t38 VSS 0.180122f
C14836 a_33496_n6659.t27 VSS 0.11863f
C14837 a_33496_n6659.n3 VSS 0.26561f
C14838 a_33496_n6659.t34 VSS 0.180122f
C14839 a_33496_n6659.t23 VSS 0.11863f
C14840 a_33496_n6659.n4 VSS 0.302075f
C14841 a_33496_n6659.t37 VSS 0.180122f
C14842 a_33496_n6659.t26 VSS 0.11863f
C14843 a_33496_n6659.n5 VSS 0.302075f
C14844 a_33496_n6659.t19 VSS 0.180122f
C14845 a_33496_n6659.t28 VSS 0.180122f
C14846 a_33496_n6659.t10 VSS 0.11863f
C14847 a_33496_n6659.n6 VSS 0.26561f
C14848 a_33496_n6659.t25 VSS 0.180122f
C14849 a_33496_n6659.t16 VSS 0.11863f
C14850 a_33496_n6659.n7 VSS 0.302075f
C14851 a_33496_n6659.t30 VSS 0.180122f
C14852 a_33496_n6659.t20 VSS 0.11863f
C14853 a_33496_n6659.n8 VSS 0.302075f
C14854 a_33496_n6659.t32 VSS 0.180122f
C14855 a_33496_n6659.t21 VSS 0.11863f
C14856 a_33496_n6659.n9 VSS -0.565154f
C14857 a_33496_n6659.t39 VSS 0.180122f
C14858 a_33496_n6659.t17 VSS 0.11863f
C14859 a_33496_n6659.n10 VSS 0.302075f
C14860 a_33496_n6659.t12 VSS 0.180122f
C14861 a_33496_n6659.t35 VSS 0.11863f
C14862 a_33496_n6659.n11 VSS 0.302075f
C14863 a_33496_n6659.t8 VSS 0.180122f
C14864 a_33496_n6659.t29 VSS 0.11863f
C14865 a_33496_n6659.n12 VSS 0.302075f
C14866 a_33496_n6659.t9 VSS 0.180122f
C14867 a_33496_n6659.t31 VSS 0.11863f
C14868 a_33496_n6659.n13 VSS 0.302075f
C14869 a_33496_n6659.t22 VSS 0.180122f
C14870 a_33496_n6659.t36 VSS 0.11863f
C14871 a_33496_n6659.n14 VSS 0.302075f
C14872 a_33496_n6659.t18 VSS 0.180122f
C14873 a_33496_n6659.t11 VSS 0.11863f
C14874 a_33496_n6659.n15 VSS 0.302075f
C14875 a_33496_n6659.t24 VSS 0.180122f
C14876 a_33496_n6659.t15 VSS 0.118046f
C14877 a_33496_n6659.t13 VSS 0.118046f
C14878 a_33496_n6659.t33 VSS 0.180122f
C14879 a_33496_n6659.t14 VSS 0.11863f
C14880 a_26553_377.t0 VSS 0.060479f
C14881 a_26553_377.t2 VSS 0.070849f
C14882 a_26553_377.t4 VSS 0.045117f
C14883 a_26553_377.n0 VSS 1.1532f
C14884 a_26553_377.t3 VSS 0.044033f
C14885 a_26553_377.t5 VSS 0.089119f
C14886 a_26553_377.n1 VSS 0.242135f
C14887 a_26553_377.n2 VSS 2.96454f
C14888 a_26553_377.n3 VSS 0.544745f
C14889 a_26553_377.t1 VSS 0.085779f
C14890 a_38256_1564.n0 VSS 0.71669f
C14891 a_38256_1564.t4 VSS 0.036741f
C14892 a_38256_1564.t6 VSS 0.050872f
C14893 a_38256_1564.t5 VSS 0.036741f
C14894 a_38256_1564.n1 VSS 0.088469f
C14895 a_38256_1564.t3 VSS 0.024695f
C14896 a_38256_1564.t2 VSS 0.024695f
C14897 a_38256_1564.n2 VSS 0.049532f
C14898 a_38256_1564.t0 VSS 0.024695f
C14899 a_38256_1564.t1 VSS 0.024695f
C14900 a_38256_1564.n3 VSS 0.05965f
C14901 a_38256_1564.t17 VSS 0.108539f
C14902 a_38256_1564.t12 VSS 0.103204f
C14903 a_38256_1564.n4 VSS 0.168431f
C14904 a_38256_1564.t20 VSS 0.108539f
C14905 a_38256_1564.t15 VSS 0.103204f
C14906 a_38256_1564.n5 VSS -0.065636f
C14907 a_38256_1564.t23 VSS 0.108539f
C14908 a_38256_1564.t19 VSS 0.103204f
C14909 a_38256_1564.n6 VSS 0.190115f
C14910 a_38256_1564.t11 VSS 0.108539f
C14911 a_38256_1564.t9 VSS 0.103204f
C14912 a_38256_1564.n7 VSS 0.190115f
C14913 a_38256_1564.t14 VSS 0.108539f
C14914 a_38256_1564.t10 VSS 0.103204f
C14915 a_38256_1564.n8 VSS 0.190115f
C14916 a_38256_1564.t18 VSS 0.108539f
C14917 a_38256_1564.t13 VSS 0.103204f
C14918 a_38256_1564.n9 VSS 0.190115f
C14919 a_38256_1564.t8 VSS 0.108539f
C14920 a_38256_1564.t21 VSS 0.103204f
C14921 a_38256_1564.n10 VSS 0.168431f
C14922 a_38256_1564.t22 VSS 0.108539f
C14923 a_38256_1564.t16 VSS 0.103204f
C14924 a_38256_1564.n11 VSS 0.273437f
C14925 a_38256_1564.n12 VSS 0.112589f
C14926 a_38256_1564.t7 VSS 0.050872f
C14927 a_11023_n22908.n0 VSS 0.016468f
C14928 a_11023_n22908.n1 VSS 0.640198f
C14929 a_11023_n22908.n2 VSS 0.056878f
C14930 a_11023_n22908.n3 VSS 0.016571f
C14931 a_11023_n22908.n4 VSS 0.056671f
C14932 a_11023_n22908.n5 VSS 0.056464f
C14933 a_11023_n22908.n6 VSS 0.056257f
C14934 a_11023_n22908.n7 VSS 0.315152f
C14935 a_11023_n22908.n8 VSS 0.315152f
C14936 a_11023_n22908.n9 VSS 0.315152f
C14937 a_11023_n22908.n10 VSS 0.436195f
C14938 a_11023_n22908.n11 VSS 0.106969f
C14939 a_11023_n22908.n12 VSS 0.052321f
C14940 a_11023_n22908.n13 VSS 0.021957f
C14941 a_11023_n22908.n14 VSS 0.052114f
C14942 a_11023_n22908.n15 VSS 0.021957f
C14943 a_11023_n22908.n16 VSS 0.051907f
C14944 a_11023_n22908.n17 VSS 0.0517f
C14945 a_11023_n22908.t12 VSS 0.0377f
C14946 a_11023_n22908.t17 VSS 0.0377f
C14947 a_11023_n22908.t11 VSS 0.0377f
C14948 a_11023_n22908.n18 VSS 0.196436f
C14949 a_11023_n22908.t15 VSS 0.0377f
C14950 a_11023_n22908.t18 VSS 0.0377f
C14951 a_11023_n22908.n19 VSS 0.181424f
C14952 a_11023_n22908.n20 VSS 0.503298f
C14953 a_11023_n22908.t38 VSS 0.064188f
C14954 a_11023_n22908.n21 VSS 0.144341f
C14955 a_11023_n22908.t20 VSS 0.064062f
C14956 a_11023_n22908.n22 VSS 0.055918f
C14957 a_11023_n22908.t34 VSS 0.064062f
C14958 a_11023_n22908.n23 VSS 0.016571f
C14959 a_11023_n22908.n24 VSS 0.119271f
C14960 a_11023_n22908.n25 VSS 0.021957f
C14961 a_11023_n22908.n26 VSS 0.021957f
C14962 a_11023_n22908.t28 VSS 0.064062f
C14963 a_11023_n22908.t39 VSS 0.064062f
C14964 a_11023_n22908.t25 VSS 0.064062f
C14965 a_11023_n22908.t23 VSS 0.064062f
C14966 a_11023_n22908.t27 VSS 0.06392f
C14967 a_11023_n22908.t36 VSS 0.063818f
C14968 a_11023_n22908.t22 VSS 0.063818f
C14969 a_11023_n22908.t29 VSS 0.063818f
C14970 a_11023_n22908.t37 VSS 0.063818f
C14971 a_11023_n22908.t24 VSS 0.063818f
C14972 a_11023_n22908.t31 VSS 0.063818f
C14973 a_11023_n22908.t26 VSS 0.063818f
C14974 a_11023_n22908.t33 VSS 0.063818f
C14975 a_11023_n22908.t21 VSS 0.063818f
C14976 a_11023_n22908.n27 VSS 0.221496f
C14977 a_11023_n22908.t35 VSS 0.064062f
C14978 a_11023_n22908.n28 VSS 0.071939f
C14979 a_11023_n22908.n29 VSS 0.021957f
C14980 a_11023_n22908.n30 VSS 0.016571f
C14981 a_11023_n22908.t30 VSS 0.064062f
C14982 a_11023_n22908.n31 VSS 0.021957f
C14983 a_11023_n22908.n32 VSS 0.021957f
C14984 a_11023_n22908.n33 VSS 0.016571f
C14985 a_11023_n22908.t32 VSS 0.064062f
C14986 a_11023_n22908.t0 VSS 0.0377f
C14987 a_11023_n22908.t4 VSS 0.0377f
C14988 a_11023_n22908.n34 VSS 0.179009f
C14989 a_11023_n22908.t3 VSS 0.0377f
C14990 a_11023_n22908.t6 VSS 0.0377f
C14991 a_11023_n22908.n35 VSS 0.179009f
C14992 a_11023_n22908.t2 VSS 0.0377f
C14993 a_11023_n22908.t9 VSS 0.0377f
C14994 a_11023_n22908.n36 VSS 0.179009f
C14995 a_11023_n22908.t5 VSS 0.0377f
C14996 a_11023_n22908.t8 VSS 0.0377f
C14997 a_11023_n22908.n37 VSS 0.179009f
C14998 a_11023_n22908.t7 VSS 0.0377f
C14999 a_11023_n22908.t1 VSS 0.0377f
C15000 a_11023_n22908.n38 VSS 0.198821f
C15001 a_11023_n22908.n39 VSS 0.696191f
C15002 a_11023_n22908.n40 VSS 0.29804f
C15003 a_11023_n22908.n41 VSS 0.29804f
C15004 a_11023_n22908.n42 VSS 0.414463f
C15005 a_11023_n22908.n43 VSS 0.718664f
C15006 a_11023_n22908.t10 VSS 0.0377f
C15007 a_11023_n22908.t14 VSS 0.0377f
C15008 a_11023_n22908.n44 VSS 0.181424f
C15009 a_11023_n22908.n45 VSS 0.319464f
C15010 a_11023_n22908.t13 VSS 0.0377f
C15011 a_11023_n22908.t16 VSS 0.0377f
C15012 a_11023_n22908.n46 VSS 0.181424f
C15013 a_11023_n22908.n47 VSS 0.184638f
C15014 a_11023_n22908.n48 VSS 0.184636f
C15015 a_11023_n22908.n49 VSS 0.181426f
C15016 a_11023_n22908.t19 VSS 0.0377f
C15017 a_13623_n22908.n0 VSS 6.32574f
C15018 a_13623_n22908.t5 VSS 0.02658f
C15019 a_13623_n22908.t7 VSS 0.029274f
C15020 a_13623_n22908.t4 VSS 0.029221f
C15021 a_13623_n22908.t6 VSS 0.02658f
C15022 a_13623_n22908.t3 VSS 0.037756f
C15023 a_13623_n22908.n1 VSS 4.5713f
C15024 a_13623_n22908.t0 VSS 0.036004f
C15025 a_13623_n22908.t2 VSS 0.03277f
C15026 a_13623_n22908.t1 VSS 0.03277f
C15027 a_13623_n22908.t14 VSS 0.038344f
C15028 a_13623_n22908.t17 VSS 0.03849f
C15029 a_13623_n22908.t30 VSS 0.038344f
C15030 a_13623_n22908.t35 VSS 0.03849f
C15031 a_13623_n22908.t20 VSS 0.038344f
C15032 a_13623_n22908.t24 VSS 0.03849f
C15033 a_13623_n22908.t9 VSS 0.038344f
C15034 a_13623_n22908.t13 VSS 0.03849f
C15035 a_13623_n22908.t29 VSS 0.038344f
C15036 a_13623_n22908.t33 VSS 0.03849f
C15037 a_13623_n22908.t8 VSS 0.038344f
C15038 a_13623_n22908.t22 VSS 0.038344f
C15039 a_13623_n22908.t15 VSS 0.038344f
C15040 a_13623_n22908.t31 VSS 0.038344f
C15041 a_13623_n22908.t25 VSS 0.038562f
C15042 a_13623_n22908.t27 VSS 0.038483f
C15043 a_13623_n22908.t10 VSS 0.038344f
C15044 a_13623_n22908.t19 VSS 0.038344f
C15045 a_13623_n22908.t12 VSS 0.038344f
C15046 a_13623_n22908.t23 VSS 0.038344f
C15047 a_13623_n22908.t34 VSS 0.038344f
C15048 a_13623_n22908.t16 VSS 0.038344f
C15049 a_13623_n22908.t26 VSS 0.038344f
C15050 a_13623_n22908.t37 VSS 0.038344f
C15051 a_13623_n22908.t32 VSS 0.038344f
C15052 a_13623_n22908.t21 VSS 0.038362f
C15053 a_13623_n22908.t36 VSS 0.03849f
C15054 a_13623_n22908.t18 VSS 0.03849f
C15055 a_13623_n22908.t28 VSS 0.03849f
C15056 a_13623_n22908.t11 VSS 0.03849f
C15057 a_13501_n9138.n0 VSS 2.0189f
C15058 a_13501_n9138.n1 VSS 3.79312f
C15059 a_13501_n9138.t12 VSS 0.041646f
C15060 a_13501_n9138.t1 VSS 0.33153f
C15061 a_13501_n9138.t13 VSS 0.321965f
C15062 a_13501_n9138.t11 VSS 0.041646f
C15063 a_13501_n9138.t15 VSS 0.041646f
C15064 a_13501_n9138.n2 VSS 0.229216f
C15065 a_13501_n9138.t6 VSS 0.041646f
C15066 a_13501_n9138.t9 VSS 0.041646f
C15067 a_13501_n9138.n3 VSS 0.223712f
C15068 a_13501_n9138.t4 VSS 0.33124f
C15069 a_13501_n9138.t14 VSS 0.325425f
C15070 a_13501_n9138.t7 VSS 0.041646f
C15071 a_13501_n9138.t0 VSS 0.041646f
C15072 a_13501_n9138.n4 VSS 0.22387f
C15073 a_13501_n9138.t17 VSS 0.041646f
C15074 a_13501_n9138.t10 VSS 0.041646f
C15075 a_13501_n9138.n5 VSS 0.228065f
C15076 a_13501_n9138.t16 VSS 0.041646f
C15077 a_13501_n9138.t19 VSS 0.041646f
C15078 a_13501_n9138.n6 VSS 0.227874f
C15079 a_13501_n9138.t8 VSS 0.041646f
C15080 a_13501_n9138.t3 VSS 0.041646f
C15081 a_13501_n9138.n7 VSS 0.22515f
C15082 a_13501_n9138.t2 VSS 0.041646f
C15083 a_13501_n9138.t5 VSS 0.041646f
C15084 a_13501_n9138.n8 VSS 0.22515f
C15085 a_13501_n9138.n9 VSS 0.228449f
C15086 a_13501_n9138.t18 VSS 0.041646f
C15087 a_11087_n10138.n0 VSS 0.96283f
C15088 a_11087_n10138.t10 VSS 0.098051f
C15089 a_11087_n10138.t2 VSS 0.100124f
C15090 a_11087_n10138.t14 VSS 0.016994f
C15091 a_11087_n10138.t17 VSS 0.096966f
C15092 a_11087_n10138.t3 VSS 0.016994f
C15093 a_11087_n10138.n1 VSS 0.232962f
C15094 a_11087_n10138.t12 VSS 0.098051f
C15095 a_11087_n10138.t16 VSS 0.016994f
C15096 a_11087_n10138.n2 VSS 0.080482f
C15097 a_11087_n10138.t7 VSS 0.097741f
C15098 a_11087_n10138.t15 VSS 0.016994f
C15099 a_11087_n10138.n3 VSS 0.080542f
C15100 a_11087_n10138.t20 VSS 0.098825f
C15101 a_11087_n10138.t28 VSS 0.016994f
C15102 a_11087_n10138.t22 VSS 0.09645f
C15103 a_11087_n10138.t25 VSS 0.016994f
C15104 a_11087_n10138.n4 VSS 0.27506f
C15105 a_11087_n10138.t29 VSS 0.095994f
C15106 a_11087_n10138.t23 VSS 0.016994f
C15107 a_11087_n10138.n5 VSS 0.094003f
C15108 a_11087_n10138.t26 VSS 0.096859f
C15109 a_11087_n10138.t24 VSS 0.016994f
C15110 a_11087_n10138.n6 VSS 0.094876f
C15111 a_11087_n10138.t27 VSS 0.095994f
C15112 a_11087_n10138.t21 VSS 0.016994f
C15113 a_11087_n10138.n7 VSS 0.165467f
C15114 a_11087_n10138.t30 VSS 4.13039f
C15115 a_11087_n10138.t31 VSS 4.28595f
C15116 a_11087_n10138.t11 VSS 0.098262f
C15117 a_11087_n10138.t5 VSS 0.016994f
C15118 a_11087_n10138.n8 VSS 1.16718f
C15119 a_11087_n10138.t6 VSS 0.098262f
C15120 a_11087_n10138.t19 VSS 0.016994f
C15121 a_11087_n10138.n9 VSS 0.08148f
C15122 a_11087_n10138.t1 VSS 0.096869f
C15123 a_11087_n10138.t13 VSS 0.016994f
C15124 a_11087_n10138.n10 VSS 0.080758f
C15125 a_11087_n10138.t4 VSS 0.096869f
C15126 a_11087_n10138.t8 VSS 0.016994f
C15127 a_11087_n10138.n11 VSS 0.081178f
C15128 a_11087_n10138.t18 VSS 0.096869f
C15129 a_11087_n10138.t9 VSS 0.016994f
C15130 a_11087_n10138.n12 VSS 0.110057f
C15131 a_11087_n10138.n13 VSS 0.340848f
C15132 a_11087_n10138.n14 VSS 0.218849f
C15133 a_11087_n10138.t0 VSS 0.016994f
C15134 a_13623_n9518.n0 VSS 6.17664f
C15135 a_13623_n9518.t5 VSS 0.042606f
C15136 a_13623_n9518.t1 VSS 0.038755f
C15137 a_13623_n9518.t7 VSS 0.038755f
C15138 a_13623_n9518.t0 VSS 0.042682f
C15139 a_13623_n9518.t6 VSS 0.05505f
C15140 a_13623_n9518.n1 VSS 3.27166f
C15141 a_13623_n9518.t2 VSS 0.050864f
C15142 a_13623_n9518.t4 VSS 0.04778f
C15143 a_13623_n9518.t3 VSS 0.055529f
C15144 a_13623_n9518.t10 VSS 0.055907f
C15145 a_13623_n9518.t24 VSS 0.056121f
C15146 a_13623_n9518.t26 VSS 0.055907f
C15147 a_13623_n9518.t12 VSS 0.056121f
C15148 a_13623_n9518.t17 VSS 0.055907f
C15149 a_13623_n9518.t16 VSS 0.056121f
C15150 a_13623_n9518.t34 VSS 0.055907f
C15151 a_13623_n9518.t25 VSS 0.055907f
C15152 a_13623_n9518.t32 VSS 0.055907f
C15153 a_13623_n9518.t19 VSS 0.055907f
C15154 a_13623_n9518.t11 VSS 0.055907f
C15155 a_13623_n9518.t27 VSS 0.055907f
C15156 a_13623_n9518.t36 VSS 0.056225f
C15157 a_13623_n9518.t23 VSS 0.05611f
C15158 a_13623_n9518.t35 VSS 0.055907f
C15159 a_13623_n9518.t15 VSS 0.055907f
C15160 a_13623_n9518.t8 VSS 0.055907f
C15161 a_13623_n9518.t21 VSS 0.055907f
C15162 a_13623_n9518.t30 VSS 0.055907f
C15163 a_13623_n9518.t13 VSS 0.055907f
C15164 a_13623_n9518.t22 VSS 0.055907f
C15165 a_13623_n9518.t31 VSS 0.055907f
C15166 a_13623_n9518.t28 VSS 0.055907f
C15167 a_13623_n9518.t18 VSS 0.055934f
C15168 a_13623_n9518.t29 VSS 0.056121f
C15169 a_13623_n9518.t14 VSS 0.056121f
C15170 a_13623_n9518.t37 VSS 0.056121f
C15171 a_13623_n9518.t20 VSS 0.056121f
C15172 a_13623_n9518.t9 VSS 0.056121f
C15173 a_13623_n9518.t33 VSS 0.056121f
C15174 OUT[5].t4 VSS 0.016573f
C15175 OUT[5].t3 VSS 0.016573f
C15176 OUT[5].n0 VSS 0.033261f
C15177 OUT[5].t2 VSS 0.016573f
C15178 OUT[5].t0 VSS 0.016573f
C15179 OUT[5].n1 VSS 0.033261f
C15180 OUT[5].t7 VSS 0.016573f
C15181 OUT[5].t6 VSS 0.016573f
C15182 OUT[5].n2 VSS 0.039859f
C15183 OUT[5].n3 VSS 0.182038f
C15184 OUT[5].t14 VSS 0.034141f
C15185 OUT[5].t13 VSS 0.024657f
C15186 OUT[5].n4 VSS 0.059536f
C15187 OUT[5].t11 VSS 0.024657f
C15188 OUT[5].t15 VSS 0.034141f
C15189 OUT[5].n5 VSS 0.074254f
C15190 OUT[5].n6 VSS 0.186805f
C15191 OUT[5].t12 VSS 0.034141f
C15192 OUT[5].t10 VSS 0.024657f
C15193 OUT[5].n7 VSS 0.059536f
C15194 OUT[5].t9 VSS 0.034141f
C15195 OUT[5].t8 VSS 0.024657f
C15196 OUT[5].n8 VSS 0.075313f
C15197 OUT[5].n9 VSS 0.190471f
C15198 OUT[5].n10 VSS 0.14639f
C15199 OUT[5].n11 VSS 0.14639f
C15200 OUT[5].n12 VSS 0.104419f
C15201 OUT[5].t1 VSS 0.016573f
C15202 OUT[5].t5 VSS 0.016573f
C15203 OUT[5].n13 VSS 0.033146f
C15204 OUT[5].n14 VSS 0.311395f
C15205 a_44640_1944.n0 VSS 0.733362f
C15206 a_44640_1944.t4 VSS 0.052055f
C15207 a_44640_1944.t0 VSS 0.025269f
C15208 a_44640_1944.t3 VSS 0.025269f
C15209 a_44640_1944.n1 VSS 0.050683f
C15210 a_44640_1944.t2 VSS 0.025269f
C15211 a_44640_1944.t1 VSS 0.025269f
C15212 a_44640_1944.n2 VSS 0.061037f
C15213 a_44640_1944.t8 VSS 0.105604f
C15214 a_44640_1944.t16 VSS 0.111063f
C15215 a_44640_1944.n3 VSS 0.172348f
C15216 a_44640_1944.t9 VSS 0.105604f
C15217 a_44640_1944.t17 VSS 0.111063f
C15218 a_44640_1944.n4 VSS -0.067162f
C15219 a_44640_1944.t21 VSS 0.105604f
C15220 a_44640_1944.t13 VSS 0.111063f
C15221 a_44640_1944.n5 VSS 0.194536f
C15222 a_44640_1944.t23 VSS 0.105604f
C15223 a_44640_1944.t15 VSS 0.111063f
C15224 a_44640_1944.n6 VSS 0.194536f
C15225 a_44640_1944.t19 VSS 0.105604f
C15226 a_44640_1944.t11 VSS 0.111063f
C15227 a_44640_1944.n7 VSS 0.194536f
C15228 a_44640_1944.t20 VSS 0.105604f
C15229 a_44640_1944.t12 VSS 0.111063f
C15230 a_44640_1944.n8 VSS 0.194536f
C15231 a_44640_1944.t18 VSS 0.105604f
C15232 a_44640_1944.t10 VSS 0.111063f
C15233 a_44640_1944.n9 VSS 0.172348f
C15234 a_44640_1944.t22 VSS 0.105604f
C15235 a_44640_1944.t14 VSS 0.111063f
C15236 a_44640_1944.n10 VSS 0.279795f
C15237 a_44640_1944.t6 VSS 0.052055f
C15238 a_44640_1944.t5 VSS 0.037595f
C15239 a_44640_1944.n11 VSS 0.115207f
C15240 a_44640_1944.n12 VSS 0.090526f
C15241 a_44640_1944.t7 VSS 0.037595f
C15242 a_10712_4516.n0 VSS 0.282683f
C15243 a_10712_4516.n1 VSS 0.312298f
C15244 a_10712_4516.n2 VSS 0.282683f
C15245 a_10712_4516.n3 VSS 0.282683f
C15246 a_10712_4516.n4 VSS 0.260649f
C15247 a_10712_4516.t21 VSS 0.034407f
C15248 a_10712_4516.t31 VSS 0.021231f
C15249 a_10712_4516.t30 VSS 0.019402f
C15250 a_10712_4516.n5 VSS 0.107257f
C15251 a_10712_4516.t49 VSS 0.024399f
C15252 a_10712_4516.t43 VSS 0.046317f
C15253 a_10712_4516.n6 VSS 0.104263f
C15254 a_10712_4516.n7 VSS 2.07384f
C15255 a_10712_4516.t26 VSS 0.034407f
C15256 a_10712_4516.t25 VSS 0.034407f
C15257 a_10712_4516.n8 VSS 0.157337f
C15258 a_10712_4516.n9 VSS 3.71419f
C15259 a_10712_4516.t23 VSS 0.034407f
C15260 a_10712_4516.t22 VSS 0.034407f
C15261 a_10712_4516.n10 VSS 0.157337f
C15262 a_10712_4516.n11 VSS 0.107293f
C15263 a_10712_4516.t20 VSS 0.034407f
C15264 a_10712_4516.t28 VSS 0.034407f
C15265 a_10712_4516.n12 VSS 0.157337f
C15266 a_10712_4516.n13 VSS 0.107293f
C15267 a_10712_4516.t38 VSS 0.058243f
C15268 a_10712_4516.t46 VSS 0.058466f
C15269 a_10712_4516.t39 VSS 0.058243f
C15270 a_10712_4516.t37 VSS 0.058243f
C15271 a_10712_4516.t44 VSS 0.058243f
C15272 a_10712_4516.t47 VSS 0.058243f
C15273 a_10712_4516.t51 VSS 0.058243f
C15274 a_10712_4516.t53 VSS 0.058243f
C15275 a_10712_4516.t35 VSS 0.058243f
C15276 a_10712_4516.t32 VSS 0.058243f
C15277 a_10712_4516.t34 VSS 0.058243f
C15278 a_10712_4516.t41 VSS 0.058466f
C15279 a_10712_4516.t40 VSS 0.058466f
C15280 a_10712_4516.t42 VSS 0.058466f
C15281 a_10712_4516.t36 VSS 0.058466f
C15282 a_10712_4516.t33 VSS 0.058466f
C15283 a_10712_4516.t52 VSS 0.058466f
C15284 a_10712_4516.t50 VSS 0.058466f
C15285 a_10712_4516.t45 VSS 0.058466f
C15286 a_10712_4516.t48 VSS 0.058466f
C15287 a_10712_4516.t7 VSS 0.034407f
C15288 a_10712_4516.t0 VSS 0.034407f
C15289 a_10712_4516.n14 VSS 0.185113f
C15290 a_10712_4516.t3 VSS 0.034407f
C15291 a_10712_4516.t5 VSS 0.034407f
C15292 a_10712_4516.n15 VSS 0.185113f
C15293 a_10712_4516.t4 VSS 0.034407f
C15294 a_10712_4516.t6 VSS 0.034407f
C15295 a_10712_4516.n16 VSS 0.185113f
C15296 a_10712_4516.t1 VSS 0.034407f
C15297 a_10712_4516.t2 VSS 0.034407f
C15298 a_10712_4516.n17 VSS 0.185113f
C15299 a_10712_4516.t8 VSS 0.034407f
C15300 a_10712_4516.t9 VSS 0.034407f
C15301 a_10712_4516.n18 VSS 0.185113f
C15302 a_10712_4516.t18 VSS 0.034407f
C15303 a_10712_4516.t17 VSS 0.034407f
C15304 a_10712_4516.n19 VSS 0.154043f
C15305 a_10712_4516.n20 VSS 0.34581f
C15306 a_10712_4516.t15 VSS 0.034407f
C15307 a_10712_4516.t14 VSS 0.034407f
C15308 a_10712_4516.n21 VSS 0.154043f
C15309 a_10712_4516.n22 VSS 0.349164f
C15310 a_10712_4516.t12 VSS 0.034407f
C15311 a_10712_4516.t10 VSS 0.034407f
C15312 a_10712_4516.n23 VSS 0.154043f
C15313 a_10712_4516.n24 VSS 0.349164f
C15314 a_10712_4516.t13 VSS 0.034407f
C15315 a_10712_4516.t11 VSS 0.034407f
C15316 a_10712_4516.n25 VSS 0.154043f
C15317 a_10712_4516.n26 VSS 0.349164f
C15318 a_10712_4516.t19 VSS 0.034407f
C15319 a_10712_4516.t16 VSS 0.034407f
C15320 a_10712_4516.n27 VSS 0.154043f
C15321 a_10712_4516.n28 VSS 0.379287f
C15322 a_10712_4516.n29 VSS 0.43096f
C15323 a_10712_4516.t27 VSS 0.034407f
C15324 a_10712_4516.t24 VSS 0.034407f
C15325 a_10712_4516.n30 VSS 0.157337f
C15326 a_10712_4516.n31 VSS 0.160925f
C15327 a_10712_4516.n32 VSS 0.107293f
C15328 a_10712_4516.n33 VSS 0.157337f
C15329 a_10712_4516.t29 VSS 0.034407f
C15330 a_10778_2852.t6 VSS 0.225803f
C15331 a_10778_2852.t3 VSS 0.222606f
C15332 a_10778_2852.t7 VSS 0.222606f
C15333 a_10778_2852.t8 VSS 0.222606f
C15334 a_10778_2852.t1 VSS 0.222606f
C15335 a_10778_2852.t0 VSS 0.219917f
C15336 a_10778_2852.t14 VSS 0.242144f
C15337 a_10778_2852.t2 VSS 0.219917f
C15338 a_10778_2852.t13 VSS 0.242144f
C15339 a_10778_2852.t9 VSS 0.219917f
C15340 a_10778_2852.t12 VSS 0.242144f
C15341 a_10778_2852.t4 VSS 0.219917f
C15342 a_10778_2852.t10 VSS 0.242144f
C15343 a_10778_2852.t5 VSS 0.219917f
C15344 a_10778_2852.t11 VSS 0.242144f
C15345 a_10778_2852.n0 VSS 1.27813f
C15346 a_10778_2852.n1 VSS 1.46912f
C15347 a_10778_2852.n2 VSS 0.875998f
C15348 a_10778_2852.n3 VSS 0.709168f
C15349 a_10778_2852.t16 VSS 0.051953f
C15350 a_10778_2852.t22 VSS 0.052152f
C15351 a_10778_2852.t17 VSS 0.051953f
C15352 a_10778_2852.t24 VSS 0.052152f
C15353 a_10778_2852.t23 VSS 0.051953f
C15354 a_10778_2852.t27 VSS 0.052152f
C15355 a_10778_2852.t25 VSS 0.051953f
C15356 a_10778_2852.t30 VSS 0.052152f
C15357 a_10778_2852.t29 VSS 0.051953f
C15358 a_10778_2852.t34 VSS 0.052152f
C15359 a_10778_2852.t33 VSS 0.051953f
C15360 a_10778_2852.t19 VSS 0.052152f
C15361 a_10778_2852.t28 VSS 0.051953f
C15362 a_10778_2852.t32 VSS 0.052152f
C15363 a_10778_2852.t31 VSS 0.051953f
C15364 a_10778_2852.t18 VSS 0.052152f
C15365 a_10778_2852.t15 VSS 0.051953f
C15366 a_10778_2852.t21 VSS 0.052152f
C15367 a_10778_2852.t20 VSS 0.051953f
C15368 a_10778_2852.t26 VSS 0.052152f
C15369 a_26388_n17606.t1 VSS 0.626206f
C15370 a_26388_n17606.n0 VSS 0.038283f
C15371 a_26388_n17606.n1 VSS 0.510238f
C15372 a_26388_n17606.t0 VSS 0.01045f
C15373 a_26388_n17606.t5 VSS 0.024337f
C15374 a_26388_n17606.t7 VSS 0.022646f
C15375 a_26388_n17606.n2 VSS 0.098809f
C15376 a_26388_n17606.t9 VSS 0.013935f
C15377 a_26388_n17606.t6 VSS 0.012735f
C15378 a_26388_n17606.t4 VSS 0.012735f
C15379 a_26388_n17606.t13 VSS 0.013935f
C15380 a_26388_n17606.n3 VSS 0.079608f
C15381 a_26388_n17606.t3 VSS 0.025965f
C15382 a_26388_n17606.t10 VSS 0.030472f
C15383 a_26388_n17606.n4 VSS 0.049615f
C15384 a_26388_n17606.n5 VSS 0.302206f
C15385 a_26388_n17606.t12 VSS 0.014204f
C15386 a_26388_n17606.t2 VSS 0.012731f
C15387 a_26388_n17606.n6 VSS 0.035653f
C15388 a_26388_n17606.n7 VSS 0.21629f
C15389 a_26388_n17606.t8 VSS 0.028948f
C15390 a_26388_n17606.t11 VSS 0.026244f
C15391 a_26388_n17606.n8 VSS 0.054511f
C15392 a_26388_n17606.n9 VSS 0.739243f
C15393 a_11087_n18172.n0 VSS 0.57197f
C15394 a_11087_n18172.n1 VSS 0.571772f
C15395 a_11087_n18172.t26 VSS 0.014027f
C15396 a_11087_n18172.t17 VSS 0.014027f
C15397 a_11087_n18172.t15 VSS 0.014027f
C15398 a_11087_n18172.n2 VSS 0.068614f
C15399 a_11087_n18172.t19 VSS 0.014027f
C15400 a_11087_n18172.t12 VSS 0.014027f
C15401 a_11087_n18172.n3 VSS 0.066007f
C15402 a_11087_n18172.n4 VSS 0.192283f
C15403 a_11087_n18172.t16 VSS 0.014027f
C15404 a_11087_n18172.t10 VSS 0.014027f
C15405 a_11087_n18172.n5 VSS 0.066903f
C15406 a_11087_n18172.n6 VSS 0.066428f
C15407 a_11087_n18172.t13 VSS 0.014027f
C15408 a_11087_n18172.t11 VSS 0.014027f
C15409 a_11087_n18172.n7 VSS 0.066647f
C15410 a_11087_n18172.n8 VSS 0.066478f
C15411 a_11087_n18172.t14 VSS 0.014027f
C15412 a_11087_n18172.t18 VSS 0.014027f
C15413 a_11087_n18172.n9 VSS 0.066903f
C15414 a_11087_n18172.n10 VSS 0.180634f
C15415 a_11087_n18172.t9 VSS 0.014027f
C15416 a_11087_n18172.t7 VSS 0.014027f
C15417 a_11087_n18172.n11 VSS 0.067542f
C15418 a_11087_n18172.t1 VSS 0.014027f
C15419 a_11087_n18172.t4 VSS 0.014027f
C15420 a_11087_n18172.n12 VSS 0.065582f
C15421 a_11087_n18172.n13 VSS 0.22703f
C15422 a_11087_n18172.t8 VSS 0.014027f
C15423 a_11087_n18172.t2 VSS 0.014027f
C15424 a_11087_n18172.n14 VSS 0.065205f
C15425 a_11087_n18172.n15 VSS 0.077588f
C15426 a_11087_n18172.t5 VSS 0.014027f
C15427 a_11087_n18172.t3 VSS 0.014027f
C15428 a_11087_n18172.n16 VSS 0.065919f
C15429 a_11087_n18172.n17 VSS 0.078309f
C15430 a_11087_n18172.t6 VSS 0.014027f
C15431 a_11087_n18172.t0 VSS 0.014027f
C15432 a_11087_n18172.n18 VSS 0.065205f
C15433 a_11087_n18172.n19 VSS 0.136734f
C15434 a_11087_n18172.n20 VSS 0.281171f
C15435 a_11087_n18172.t35 VSS 3.68956f
C15436 a_11087_n18172.t33 VSS 3.57447f
C15437 a_11087_n18172.n21 VSS 0.715158f
C15438 a_11087_n18172.t32 VSS 3.54024f
C15439 a_11087_n18172.t36 VSS 3.69935f
C15440 a_11087_n18172.n22 VSS 1.00626f
C15441 a_11087_n18172.t37 VSS 4.04337f
C15442 a_11087_n18172.t34 VSS 3.49998f
C15443 a_11087_n18172.n23 VSS 0.73941f
C15444 a_11087_n18172.t30 VSS 3.53756f
C15445 a_11087_n18172.t31 VSS 3.49937f
C15446 a_11087_n18172.n24 VSS 0.633447f
C15447 a_11087_n18172.n25 VSS 0.908383f
C15448 a_11087_n18172.t28 VSS 0.014027f
C15449 a_11087_n18172.t22 VSS 0.014027f
C15450 a_11087_n18172.n26 VSS 0.067077f
C15451 a_11087_n18172.n27 VSS 0.354035f
C15452 a_11087_n18172.t21 VSS 0.014027f
C15453 a_11087_n18172.t25 VSS 0.014027f
C15454 a_11087_n18172.n28 VSS 0.067077f
C15455 a_11087_n18172.n29 VSS 0.067252f
C15456 a_11087_n18172.t24 VSS 0.014027f
C15457 a_11087_n18172.t27 VSS 0.014027f
C15458 a_11087_n18172.n30 VSS 0.065927f
C15459 a_11087_n18172.n31 VSS 0.066656f
C15460 a_11087_n18172.t23 VSS 0.014027f
C15461 a_11087_n18172.t20 VSS 0.014027f
C15462 a_11087_n18172.n32 VSS 0.065927f
C15463 a_11087_n18172.n33 VSS 0.067003f
C15464 a_11087_n18172.n34 VSS 0.090839f
C15465 a_11087_n18172.n35 VSS 0.065927f
C15466 a_11087_n18172.t29 VSS 0.014027f
C15467 a_11023_n17552.n0 VSS 0.016166f
C15468 a_11023_n17552.n1 VSS 0.628451f
C15469 a_11023_n17552.n2 VSS 0.055834f
C15470 a_11023_n17552.n3 VSS 0.016267f
C15471 a_11023_n17552.n4 VSS 0.055631f
C15472 a_11023_n17552.n5 VSS 0.055428f
C15473 a_11023_n17552.n6 VSS 0.055225f
C15474 a_11023_n17552.n7 VSS 0.309369f
C15475 a_11023_n17552.n8 VSS 0.309369f
C15476 a_11023_n17552.n9 VSS 0.309369f
C15477 a_11023_n17552.n10 VSS 0.428191f
C15478 a_11023_n17552.n11 VSS 0.105007f
C15479 a_11023_n17552.n12 VSS 0.051361f
C15480 a_11023_n17552.n13 VSS 0.021554f
C15481 a_11023_n17552.n14 VSS 0.051158f
C15482 a_11023_n17552.n15 VSS 0.021554f
C15483 a_11023_n17552.n16 VSS 0.050954f
C15484 a_11023_n17552.n17 VSS 0.050751f
C15485 a_11023_n17552.t16 VSS 0.037008f
C15486 a_11023_n17552.t14 VSS 0.037008f
C15487 a_11023_n17552.t18 VSS 0.037008f
C15488 a_11023_n17552.n18 VSS 0.192832f
C15489 a_11023_n17552.t12 VSS 0.037008f
C15490 a_11023_n17552.t15 VSS 0.037008f
C15491 a_11023_n17552.n19 VSS 0.178095f
C15492 a_11023_n17552.n20 VSS 0.494064f
C15493 a_11023_n17552.t25 VSS 0.06301f
C15494 a_11023_n17552.n21 VSS 0.141693f
C15495 a_11023_n17552.t27 VSS 0.062887f
C15496 a_11023_n17552.n22 VSS 0.054892f
C15497 a_11023_n17552.t21 VSS 0.062887f
C15498 a_11023_n17552.n23 VSS 0.016267f
C15499 a_11023_n17552.n24 VSS 0.117082f
C15500 a_11023_n17552.n25 VSS 0.021554f
C15501 a_11023_n17552.n26 VSS 0.021554f
C15502 a_11023_n17552.t35 VSS 0.062887f
C15503 a_11023_n17552.t26 VSS 0.062887f
C15504 a_11023_n17552.t32 VSS 0.062887f
C15505 a_11023_n17552.t30 VSS 0.062887f
C15506 a_11023_n17552.t34 VSS 0.062747f
C15507 a_11023_n17552.t23 VSS 0.062647f
C15508 a_11023_n17552.t29 VSS 0.062647f
C15509 a_11023_n17552.t36 VSS 0.062647f
C15510 a_11023_n17552.t24 VSS 0.062647f
C15511 a_11023_n17552.t31 VSS 0.062647f
C15512 a_11023_n17552.t38 VSS 0.062647f
C15513 a_11023_n17552.t33 VSS 0.062647f
C15514 a_11023_n17552.t20 VSS 0.062647f
C15515 a_11023_n17552.t28 VSS 0.062647f
C15516 a_11023_n17552.n27 VSS 0.217432f
C15517 a_11023_n17552.t22 VSS 0.062887f
C15518 a_11023_n17552.n28 VSS 0.070619f
C15519 a_11023_n17552.n29 VSS 0.021554f
C15520 a_11023_n17552.n30 VSS 0.016267f
C15521 a_11023_n17552.t37 VSS 0.062887f
C15522 a_11023_n17552.n31 VSS 0.021554f
C15523 a_11023_n17552.n32 VSS 0.021554f
C15524 a_11023_n17552.n33 VSS 0.016267f
C15525 a_11023_n17552.t39 VSS 0.062887f
C15526 a_11023_n17552.t7 VSS 0.037008f
C15527 a_11023_n17552.t1 VSS 0.037008f
C15528 a_11023_n17552.n34 VSS 0.175725f
C15529 a_11023_n17552.t0 VSS 0.037008f
C15530 a_11023_n17552.t3 VSS 0.037008f
C15531 a_11023_n17552.n35 VSS 0.175725f
C15532 a_11023_n17552.t9 VSS 0.037008f
C15533 a_11023_n17552.t6 VSS 0.037008f
C15534 a_11023_n17552.n36 VSS 0.175725f
C15535 a_11023_n17552.t2 VSS 0.037008f
C15536 a_11023_n17552.t5 VSS 0.037008f
C15537 a_11023_n17552.n37 VSS 0.175725f
C15538 a_11023_n17552.t4 VSS 0.037008f
C15539 a_11023_n17552.t8 VSS 0.037008f
C15540 a_11023_n17552.n38 VSS 0.195173f
C15541 a_11023_n17552.n39 VSS 0.683417f
C15542 a_11023_n17552.n40 VSS 0.292571f
C15543 a_11023_n17552.n41 VSS 0.292571f
C15544 a_11023_n17552.n42 VSS 0.406859f
C15545 a_11023_n17552.n43 VSS 0.705478f
C15546 a_11023_n17552.t17 VSS 0.037008f
C15547 a_11023_n17552.t11 VSS 0.037008f
C15548 a_11023_n17552.n44 VSS 0.178095f
C15549 a_11023_n17552.n45 VSS 0.313602f
C15550 a_11023_n17552.t10 VSS 0.037008f
C15551 a_11023_n17552.t13 VSS 0.037008f
C15552 a_11023_n17552.n46 VSS 0.178095f
C15553 a_11023_n17552.n47 VSS 0.18125f
C15554 a_11023_n17552.n48 VSS 0.181248f
C15555 a_11023_n17552.n49 VSS 0.178097f
C15556 a_11023_n17552.t19 VSS 0.037008f
C15557 a_21692_n5468.n0 VSS 0.555747f
C15558 a_21692_n5468.n1 VSS 0.28906f
C15559 a_21692_n5468.n2 VSS 0.201659f
C15560 a_21692_n5468.t12 VSS 0.041975f
C15561 a_21692_n5468.t14 VSS 0.041975f
C15562 a_21692_n5468.t10 VSS 0.041975f
C15563 a_21692_n5468.n3 VSS 0.085002f
C15564 a_21692_n5468.t11 VSS 0.041975f
C15565 a_21692_n5468.t9 VSS 0.041975f
C15566 a_21692_n5468.n4 VSS 0.0864f
C15567 a_21692_n5468.t28 VSS 0.052258f
C15568 a_21692_n5468.t20 VSS 0.061644f
C15569 a_21692_n5468.n5 VSS 0.265472f
C15570 a_21692_n5468.t29 VSS 0.06045f
C15571 a_21692_n5468.t26 VSS 0.054344f
C15572 a_21692_n5468.n6 VSS 0.128082f
C15573 a_21692_n5468.t27 VSS 0.054597f
C15574 a_21692_n5468.t31 VSS 0.060211f
C15575 a_21692_n5468.n7 VSS 0.144304f
C15576 a_21692_n5468.t32 VSS 0.06045f
C15577 a_21692_n5468.t16 VSS 0.054344f
C15578 a_21692_n5468.n8 VSS 0.126316f
C15579 a_21692_n5468.n9 VSS 0.569043f
C15580 a_21692_n5468.n10 VSS 0.608363f
C15581 a_21692_n5468.t23 VSS 0.06045f
C15582 a_21692_n5468.t19 VSS 0.054344f
C15583 a_21692_n5468.n11 VSS 0.164831f
C15584 a_21692_n5468.n12 VSS 1.37551f
C15585 a_21692_n5468.t21 VSS 0.052258f
C15586 a_21692_n5468.t17 VSS 0.061644f
C15587 a_21692_n5468.n13 VSS 0.120547f
C15588 a_21692_n5468.n14 VSS 0.729969f
C15589 a_21692_n5468.t22 VSS 0.054597f
C15590 a_21692_n5468.t30 VSS 0.060211f
C15591 a_21692_n5468.n15 VSS 0.121623f
C15592 a_21692_n5468.n16 VSS 0.85621f
C15593 a_21692_n5468.t18 VSS 0.054597f
C15594 a_21692_n5468.t25 VSS 0.060211f
C15595 a_21692_n5468.n17 VSS 0.121366f
C15596 a_21692_n5468.n18 VSS 0.720147f
C15597 a_21692_n5468.t24 VSS 0.054597f
C15598 a_21692_n5468.t33 VSS 0.060211f
C15599 a_21692_n5468.n19 VSS 0.121623f
C15600 a_21692_n5468.n20 VSS 1.1183f
C15601 a_21692_n5468.n21 VSS 1.64319f
C15602 a_21692_n5468.t2 VSS 0.010685f
C15603 a_21692_n5468.t3 VSS 0.010685f
C15604 a_21692_n5468.n22 VSS 0.021702f
C15605 a_21692_n5468.t4 VSS 0.010685f
C15606 a_21692_n5468.t5 VSS 0.010685f
C15607 a_21692_n5468.n23 VSS 0.030614f
C15608 a_21692_n5468.t1 VSS 0.010685f
C15609 a_21692_n5468.t0 VSS 0.010685f
C15610 a_21692_n5468.n24 VSS 0.021702f
C15611 a_21692_n5468.t6 VSS 0.010685f
C15612 a_21692_n5468.t7 VSS 0.010685f
C15613 a_21692_n5468.n25 VSS 0.030614f
C15614 a_21692_n5468.t8 VSS 0.041975f
C15615 a_21692_n5468.t13 VSS 0.041975f
C15616 a_21692_n5468.n26 VSS 0.104908f
C15617 a_21692_n5468.n27 VSS 0.085002f
C15618 a_21692_n5468.t15 VSS 0.041975f
C15619 a_26440_n5940.n0 VSS 0.709036f
C15620 a_26440_n5940.t3 VSS 0.042608f
C15621 a_26440_n5940.t0 VSS 0.070466f
C15622 a_26440_n5940.t1 VSS 0.079497f
C15623 a_26440_n5940.t2 VSS 0.021375f
C15624 a_26440_n5940.t8 VSS 0.04632f
C15625 a_26440_n5940.t11 VSS 0.076349f
C15626 a_26440_n5940.n1 VSS 0.111235f
C15627 a_26440_n5940.t4 VSS 0.04632f
C15628 a_26440_n5940.t14 VSS 0.076349f
C15629 a_26440_n5940.t10 VSS 0.04632f
C15630 a_26440_n5940.t7 VSS 0.076349f
C15631 a_26440_n5940.n2 VSS 0.111235f
C15632 a_26440_n5940.t12 VSS 0.04632f
C15633 a_26440_n5940.t16 VSS 0.076349f
C15634 a_26440_n5940.n3 VSS -0.029833f
C15635 a_26440_n5940.t15 VSS 0.04632f
C15636 a_26440_n5940.t9 VSS 0.076349f
C15637 a_26440_n5940.n4 VSS 0.126528f
C15638 a_26440_n5940.t17 VSS 0.04632f
C15639 a_26440_n5940.t5 VSS 0.076349f
C15640 a_26440_n5940.n5 VSS 0.126528f
C15641 a_26440_n5940.t19 VSS 0.04632f
C15642 a_26440_n5940.t13 VSS 0.076349f
C15643 a_26440_n5940.n6 VSS 0.126528f
C15644 a_26440_n5940.t18 VSS 0.04632f
C15645 a_26440_n5940.t6 VSS 0.076349f
C15646 a_26440_n5940.n7 VSS 0.12344f
C15647 a_28721_n9076.t1 VSS 0.523935f
C15648 a_28721_n9076.n0 VSS 0.581482f
C15649 a_28721_n9076.t0 VSS 0.024933f
C15650 a_28721_n9076.t6 VSS 0.079133f
C15651 a_28721_n9076.t3 VSS 0.046948f
C15652 a_28721_n9076.n1 VSS 0.33635f
C15653 a_28721_n9076.t4 VSS 0.05915f
C15654 a_28721_n9076.t7 VSS 0.080285f
C15655 a_28721_n9076.n2 VSS 0.256016f
C15656 a_28721_n9076.n3 VSS 1.36939f
C15657 a_28721_n9076.t9 VSS 0.051291f
C15658 a_28721_n9076.t5 VSS 0.08816f
C15659 a_28721_n9076.n4 VSS 0.089376f
C15660 a_28721_n9076.t8 VSS 0.053728f
C15661 a_28721_n9076.t2 VSS 0.056084f
C15662 a_28721_n9076.n5 VSS 0.103741f
C15663 a_11087_n15494.n0 VSS 1.10641f
C15664 a_11087_n15494.t23 VSS 0.0175f
C15665 a_11087_n15494.t15 VSS 0.0175f
C15666 a_11087_n15494.t13 VSS 0.0175f
C15667 a_11087_n15494.n1 VSS 0.085607f
C15668 a_11087_n15494.t17 VSS 0.0175f
C15669 a_11087_n15494.t10 VSS 0.0175f
C15670 a_11087_n15494.n2 VSS 0.082354f
C15671 a_11087_n15494.n3 VSS 0.239903f
C15672 a_11087_n15494.t14 VSS 0.0175f
C15673 a_11087_n15494.t18 VSS 0.0175f
C15674 a_11087_n15494.n4 VSS 0.083472f
C15675 a_11087_n15494.n5 VSS 0.082879f
C15676 a_11087_n15494.t11 VSS 0.0175f
C15677 a_11087_n15494.t19 VSS 0.0175f
C15678 a_11087_n15494.n6 VSS 0.083153f
C15679 a_11087_n15494.n7 VSS 0.082941f
C15680 a_11087_n15494.t12 VSS 0.0175f
C15681 a_11087_n15494.t16 VSS 0.0175f
C15682 a_11087_n15494.n8 VSS 0.083472f
C15683 a_11087_n15494.n9 VSS 0.225369f
C15684 a_11087_n15494.t3 VSS 0.0175f
C15685 a_11087_n15494.t5 VSS 0.0175f
C15686 a_11087_n15494.n10 VSS 0.084269f
C15687 a_11087_n15494.t1 VSS 0.0175f
C15688 a_11087_n15494.t8 VSS 0.0175f
C15689 a_11087_n15494.n11 VSS 0.081823f
C15690 a_11087_n15494.n12 VSS 0.283255f
C15691 a_11087_n15494.t4 VSS 0.0175f
C15692 a_11087_n15494.t0 VSS 0.0175f
C15693 a_11087_n15494.n13 VSS 0.081354f
C15694 a_11087_n15494.n14 VSS 0.096803f
C15695 a_11087_n15494.t7 VSS 0.0175f
C15696 a_11087_n15494.t9 VSS 0.0175f
C15697 a_11087_n15494.n15 VSS 0.082244f
C15698 a_11087_n15494.n16 VSS 0.097702f
C15699 a_11087_n15494.t6 VSS 0.0175f
C15700 a_11087_n15494.t2 VSS 0.0175f
C15701 a_11087_n15494.n17 VSS 0.081354f
C15702 a_11087_n15494.n18 VSS 0.170596f
C15703 a_11087_n15494.n19 VSS 0.350804f
C15704 a_11087_n15494.t24 VSS 0.0175f
C15705 a_11087_n15494.t27 VSS 0.0175f
C15706 a_11087_n15494.n20 VSS 0.082254f
C15707 a_11087_n15494.n21 VSS 0.113336f
C15708 a_11087_n15494.t21 VSS 0.0175f
C15709 a_11087_n15494.t28 VSS 0.0175f
C15710 a_11087_n15494.n22 VSS 0.082254f
C15711 a_11087_n15494.n23 VSS 0.083597f
C15712 a_11087_n15494.t22 VSS 0.0175f
C15713 a_11087_n15494.t25 VSS 0.0175f
C15714 a_11087_n15494.n24 VSS 0.082254f
C15715 a_11087_n15494.n25 VSS 0.083164f
C15716 a_11087_n15494.t33 VSS 5.37331f
C15717 a_11087_n15494.t32 VSS 4.26307f
C15718 a_11087_n15494.n26 VSS 1.67107f
C15719 a_11087_n15494.t30 VSS 4.73781f
C15720 a_11087_n15494.t31 VSS 4.41364f
C15721 a_11087_n15494.n27 VSS 1.26149f
C15722 a_11087_n15494.t26 VSS 0.0175f
C15723 a_11087_n15494.t20 VSS 0.0175f
C15724 a_11087_n15494.n28 VSS 0.083689f
C15725 a_11087_n15494.n29 VSS 0.510674f
C15726 a_11087_n15494.n30 VSS 0.083907f
C15727 a_11087_n15494.n31 VSS 0.083689f
C15728 a_11087_n15494.t29 VSS 0.0175f
C15729 a_11023_n14874.n0 VSS 0.904871f
C15730 a_11023_n14874.t29 VSS 0.065212f
C15731 a_11023_n14874.n1 VSS 0.782917f
C15732 a_11023_n14874.n2 VSS 1.64085f
C15733 a_11023_n14874.t9 VSS 0.219126f
C15734 a_11023_n14874.t13 VSS 0.234136f
C15735 a_11023_n14874.t4 VSS 0.0377f
C15736 a_11023_n14874.t17 VSS 0.219124f
C15737 a_11023_n14874.t10 VSS 0.0377f
C15738 a_11023_n14874.n3 VSS 0.503298f
C15739 a_11023_n14874.t31 VSS 0.064062f
C15740 a_11023_n14874.t25 VSS 0.064062f
C15741 a_11023_n14874.t39 VSS 0.064062f
C15742 a_11023_n14874.t30 VSS 0.064062f
C15743 a_11023_n14874.t36 VSS 0.064062f
C15744 a_11023_n14874.t34 VSS 0.064062f
C15745 a_11023_n14874.t38 VSS 0.06392f
C15746 a_11023_n14874.t27 VSS 0.063818f
C15747 a_11023_n14874.t33 VSS 0.063818f
C15748 a_11023_n14874.t20 VSS 0.063818f
C15749 a_11023_n14874.t28 VSS 0.063818f
C15750 a_11023_n14874.t35 VSS 0.063818f
C15751 a_11023_n14874.t22 VSS 0.063818f
C15752 a_11023_n14874.t37 VSS 0.063818f
C15753 a_11023_n14874.t24 VSS 0.063818f
C15754 a_11023_n14874.t32 VSS 0.063818f
C15755 a_11023_n14874.t26 VSS 0.064062f
C15756 a_11023_n14874.t21 VSS 0.064062f
C15757 a_11023_n14874.t23 VSS 0.064062f
C15758 a_11023_n14874.t8 VSS 0.216709f
C15759 a_11023_n14874.t1 VSS 0.0377f
C15760 a_11023_n14874.t2 VSS 0.216709f
C15761 a_11023_n14874.t16 VSS 0.0377f
C15762 a_11023_n14874.t6 VSS 0.216709f
C15763 a_11023_n14874.t11 VSS 0.0377f
C15764 a_11023_n14874.t0 VSS 0.216709f
C15765 a_11023_n14874.t12 VSS 0.0377f
C15766 a_11023_n14874.t15 VSS 0.236521f
C15767 a_11023_n14874.t7 VSS 0.0377f
C15768 a_11023_n14874.n4 VSS 0.696191f
C15769 a_11023_n14874.n5 VSS 0.29804f
C15770 a_11023_n14874.n6 VSS 0.29804f
C15771 a_11023_n14874.n7 VSS 0.414463f
C15772 a_11023_n14874.n8 VSS 0.801546f
C15773 a_11023_n14874.t5 VSS 0.219124f
C15774 a_11023_n14874.t18 VSS 0.0377f
C15775 a_11023_n14874.n9 VSS 0.319464f
C15776 a_11023_n14874.t19 VSS 0.219124f
C15777 a_11023_n14874.t14 VSS 0.0377f
C15778 a_11023_n14874.n10 VSS 0.184638f
C15779 a_11023_n14874.n11 VSS 0.184636f
C15780 a_11023_n14874.t3 VSS 0.0377f
C15781 a_13623_n17552.n0 VSS 3.55445f
C15782 a_13623_n17552.n1 VSS 0.400361f
C15783 a_13623_n17552.n2 VSS 0.430267f
C15784 a_13623_n17552.n3 VSS 2.46316f
C15785 a_13623_n17552.n4 VSS 0.289408f
C15786 a_13623_n17552.t13 VSS 0.010562f
C15787 a_13623_n17552.t10 VSS 0.010562f
C15788 a_13623_n17552.t12 VSS 0.014625f
C15789 a_13623_n17552.n5 VSS 0.025503f
C15790 a_13623_n17552.t11 VSS 0.014625f
C15791 a_13623_n17552.t9 VSS 0.010562f
C15792 a_13623_n17552.n6 VSS 0.031808f
C15793 a_13623_n17552.n7 VSS 0.014248f
C15794 a_13623_n17552.n8 VSS 0.017074f
C15795 a_13623_n17552.n9 VSS 0.014248f
C15796 a_13623_n17552.n10 VSS 0.017131f
C15797 a_13623_n17552.t14 VSS 0.010562f
C15798 a_13623_n17552.t8 VSS 0.014625f
C15799 a_13623_n17552.n11 VSS 0.026393f
C15800 a_13623_n17552.t31 VSS 0.041036f
C15801 a_13623_n17552.t34 VSS 0.041193f
C15802 a_13623_n17552.t17 VSS 0.041036f
C15803 a_13623_n17552.t37 VSS 0.041036f
C15804 a_13623_n17552.t26 VSS 0.041036f
C15805 a_13623_n17552.t16 VSS 0.041036f
C15806 a_13623_n17552.t25 VSS 0.041036f
C15807 a_13623_n17552.t39 VSS 0.041036f
C15808 a_13623_n17552.t32 VSS 0.041036f
C15809 a_13623_n17552.t18 VSS 0.041036f
C15810 a_13623_n17552.t42 VSS 0.04127f
C15811 a_13623_n17552.t44 VSS 0.041185f
C15812 a_13623_n17552.t27 VSS 0.041036f
C15813 a_13623_n17552.t36 VSS 0.041036f
C15814 a_13623_n17552.t29 VSS 0.041036f
C15815 a_13623_n17552.t40 VSS 0.041036f
C15816 a_13623_n17552.t21 VSS 0.041036f
C15817 a_13623_n17552.t33 VSS 0.041036f
C15818 a_13623_n17552.t43 VSS 0.041036f
C15819 a_13623_n17552.t24 VSS 0.041036f
C15820 a_13623_n17552.t19 VSS 0.041036f
C15821 a_13623_n17552.t38 VSS 0.041056f
C15822 a_13623_n17552.t23 VSS 0.041193f
C15823 a_13623_n17552.t35 VSS 0.041193f
C15824 a_13623_n17552.t45 VSS 0.041193f
C15825 a_13623_n17552.t28 VSS 0.041193f
C15826 a_13623_n17552.t20 VSS 0.041193f
C15827 a_13623_n17552.t30 VSS 0.041193f
C15828 a_13623_n17552.t41 VSS 0.041193f
C15829 a_13623_n17552.t22 VSS 0.041193f
C15830 a_13623_n17552.n12 VSS 0.025503f
C15831 a_13623_n17552.t15 VSS 0.014625f
C15832 a_21772_n8292.n0 VSS 0.38344f
C15833 a_21772_n8292.t6 VSS 0.019652f
C15834 a_21772_n8292.t5 VSS 0.019652f
C15835 a_21772_n8292.t4 VSS 0.027211f
C15836 a_21772_n8292.n1 VSS 0.047321f
C15837 a_21772_n8292.t2 VSS 0.013209f
C15838 a_21772_n8292.t3 VSS 0.013209f
C15839 a_21772_n8292.n2 VSS 0.026494f
C15840 a_21772_n8292.t0 VSS 0.013209f
C15841 a_21772_n8292.t1 VSS 0.013209f
C15842 a_21772_n8292.n3 VSS 0.031906f
C15843 a_21772_n8292.t18 VSS 0.058056f
C15844 a_21772_n8292.t12 VSS 0.055202f
C15845 a_21772_n8292.n4 VSS 0.090091f
C15846 a_21772_n8292.t23 VSS 0.058056f
C15847 a_21772_n8292.t17 VSS 0.055202f
C15848 a_21772_n8292.n5 VSS 0.090091f
C15849 a_21772_n8292.t13 VSS 0.058056f
C15850 a_21772_n8292.t21 VSS 0.055202f
C15851 a_21772_n8292.n6 VSS -0.035108f
C15852 a_21772_n8292.t11 VSS 0.058056f
C15853 a_21772_n8292.t22 VSS 0.055202f
C15854 a_21772_n8292.n7 VSS 0.101689f
C15855 a_21772_n8292.t14 VSS 0.058056f
C15856 a_21772_n8292.t8 VSS 0.055202f
C15857 a_21772_n8292.n8 VSS 0.101689f
C15858 a_21772_n8292.t16 VSS 0.058056f
C15859 a_21772_n8292.t10 VSS 0.055202f
C15860 a_21772_n8292.n9 VSS 0.101689f
C15861 a_21772_n8292.t19 VSS 0.058056f
C15862 a_21772_n8292.t9 VSS 0.055202f
C15863 a_21772_n8292.n10 VSS 0.101689f
C15864 a_21772_n8292.t20 VSS 0.058056f
C15865 a_21772_n8292.t15 VSS 0.055202f
C15866 a_21772_n8292.n11 VSS 0.146163f
C15867 a_21772_n8292.n12 VSS 0.060222f
C15868 a_21772_n8292.t7 VSS 0.027211f
C15869 a_11087_n7460.t24 VSS 0.025904f
C15870 a_11087_n7460.t3 VSS 0.025904f
C15871 a_11087_n7460.t8 VSS 0.025904f
C15872 a_11087_n7460.n0 VSS 0.124732f
C15873 a_11087_n7460.t1 VSS 0.025904f
C15874 a_11087_n7460.t4 VSS 0.025904f
C15875 a_11087_n7460.n1 VSS 0.121112f
C15876 a_11087_n7460.n2 VSS 0.419264f
C15877 a_11087_n7460.t7 VSS 0.025904f
C15878 a_11087_n7460.t0 VSS 0.025904f
C15879 a_11087_n7460.n3 VSS 0.120417f
C15880 a_11087_n7460.n4 VSS 0.143285f
C15881 a_11087_n7460.t5 VSS 0.025904f
C15882 a_11087_n7460.t9 VSS 0.025904f
C15883 a_11087_n7460.n5 VSS 0.121735f
C15884 a_11087_n7460.n6 VSS 0.144616f
C15885 a_11087_n7460.t2 VSS 0.025904f
C15886 a_11087_n7460.t6 VSS 0.025904f
C15887 a_11087_n7460.n7 VSS 0.120417f
C15888 a_11087_n7460.n8 VSS 0.252215f
C15889 a_11087_n7460.t30 VSS 5.61207f
C15890 a_11087_n7460.t12 VSS 0.025904f
C15891 a_11087_n7460.t18 VSS 0.025904f
C15892 a_11087_n7460.n9 VSS 0.123874f
C15893 a_11087_n7460.n10 VSS 1.81879f
C15894 a_11087_n7460.t17 VSS 0.025904f
C15895 a_11087_n7460.t15 VSS 0.025904f
C15896 a_11087_n7460.n11 VSS 0.123874f
C15897 a_11087_n7460.n12 VSS 0.124197f
C15898 a_11087_n7460.t14 VSS 0.025904f
C15899 a_11087_n7460.t11 VSS 0.025904f
C15900 a_11087_n7460.n13 VSS 0.12175f
C15901 a_11087_n7460.n14 VSS 0.123097f
C15902 a_11087_n7460.t13 VSS 0.025904f
C15903 a_11087_n7460.t19 VSS 0.025904f
C15904 a_11087_n7460.n15 VSS 0.12175f
C15905 a_11087_n7460.n16 VSS 0.123737f
C15906 a_11087_n7460.t10 VSS 0.025904f
C15907 a_11087_n7460.t16 VSS 0.025904f
C15908 a_11087_n7460.n17 VSS 0.12175f
C15909 a_11087_n7460.n18 VSS 0.167756f
C15910 a_11087_n7460.n19 VSS 0.519543f
C15911 a_11087_n7460.t25 VSS 0.025904f
C15912 a_11087_n7460.t21 VSS 0.025904f
C15913 a_11087_n7460.n20 VSS 0.123552f
C15914 a_11087_n7460.n21 VSS 0.333583f
C15915 a_11087_n7460.t22 VSS 0.025904f
C15916 a_11087_n7460.t28 VSS 0.025904f
C15917 a_11087_n7460.n22 VSS 0.12308f
C15918 a_11087_n7460.n23 VSS 0.122767f
C15919 a_11087_n7460.t20 VSS 0.025904f
C15920 a_11087_n7460.t27 VSS 0.025904f
C15921 a_11087_n7460.n24 VSS 0.123552f
C15922 a_11087_n7460.n25 VSS 0.122675f
C15923 a_11087_n7460.t26 VSS 0.025904f
C15924 a_11087_n7460.t23 VSS 0.025904f
C15925 a_11087_n7460.n26 VSS 0.121898f
C15926 a_11087_n7460.n27 VSS 0.355095f
C15927 a_11087_n7460.n28 VSS 0.126712f
C15928 a_11087_n7460.t29 VSS 0.025904f
C15929 a_13501_n6460.t10 VSS 0.307161f
C15930 a_13501_n6460.t8 VSS 0.308441f
C15931 a_13501_n6460.t11 VSS 0.307003f
C15932 a_13501_n6460.t6 VSS 0.308441f
C15933 a_13501_n6460.t2 VSS 0.311357f
C15934 a_13501_n6460.t0 VSS 0.311165f
C15935 a_13501_n6460.t4 VSS 0.31174f
C15936 a_13501_n6460.t1 VSS 0.312507f
C15937 a_13501_n6460.n0 VSS 5.81203f
C15938 a_13501_n6460.t9 VSS 0.33153f
C15939 a_13501_n6460.t3 VSS 0.321965f
C15940 a_13501_n6460.t7 VSS 0.33124f
C15941 a_13501_n6460.t5 VSS 0.325425f
C15942 a_11023_n6840.n0 VSS 0.904871f
C15943 a_11023_n6840.t27 VSS 0.065212f
C15944 a_11023_n6840.n1 VSS 0.782917f
C15945 a_11023_n6840.n2 VSS 1.64085f
C15946 a_11023_n6840.t14 VSS 0.234139f
C15947 a_11023_n6840.t20 VSS 0.064062f
C15948 a_11023_n6840.t24 VSS 0.064062f
C15949 a_11023_n6840.t29 VSS 0.064062f
C15950 a_11023_n6840.t38 VSS 0.064062f
C15951 a_11023_n6840.t33 VSS 0.064062f
C15952 a_11023_n6840.t25 VSS 0.064062f
C15953 a_11023_n6840.t26 VSS 0.06392f
C15954 a_11023_n6840.t35 VSS 0.063818f
C15955 a_11023_n6840.t31 VSS 0.063818f
C15956 a_11023_n6840.t28 VSS 0.063818f
C15957 a_11023_n6840.t37 VSS 0.063818f
C15958 a_11023_n6840.t32 VSS 0.063818f
C15959 a_11023_n6840.t22 VSS 0.063818f
C15960 a_11023_n6840.t34 VSS 0.063818f
C15961 a_11023_n6840.t30 VSS 0.063818f
C15962 a_11023_n6840.t39 VSS 0.063818f
C15963 a_11023_n6840.t36 VSS 0.064062f
C15964 a_11023_n6840.t21 VSS 0.064062f
C15965 a_11023_n6840.t23 VSS 0.064062f
C15966 a_11023_n6840.t17 VSS 0.216709f
C15967 a_11023_n6840.t1 VSS 0.0377f
C15968 a_11023_n6840.t2 VSS 0.216709f
C15969 a_11023_n6840.t7 VSS 0.0377f
C15970 a_11023_n6840.t4 VSS 0.216709f
C15971 a_11023_n6840.t12 VSS 0.0377f
C15972 a_11023_n6840.t10 VSS 0.216709f
C15973 a_11023_n6840.t0 VSS 0.0377f
C15974 a_11023_n6840.t16 VSS 0.236521f
C15975 a_11023_n6840.t6 VSS 0.0377f
C15976 a_11023_n6840.n3 VSS 0.696191f
C15977 a_11023_n6840.n4 VSS 0.29804f
C15978 a_11023_n6840.n5 VSS 0.29804f
C15979 a_11023_n6840.n6 VSS 0.414463f
C15980 a_11023_n6840.n7 VSS 0.801546f
C15981 a_11023_n6840.t5 VSS 0.219124f
C15982 a_11023_n6840.t9 VSS 0.0377f
C15983 a_11023_n6840.n8 VSS 0.319464f
C15984 a_11023_n6840.t11 VSS 0.219124f
C15985 a_11023_n6840.t15 VSS 0.0377f
C15986 a_11023_n6840.n9 VSS 0.184638f
C15987 a_11023_n6840.t13 VSS 0.219124f
C15988 a_11023_n6840.t19 VSS 0.0377f
C15989 a_11023_n6840.n10 VSS 0.184638f
C15990 a_11023_n6840.t18 VSS 0.219124f
C15991 a_11023_n6840.t8 VSS 0.0377f
C15992 a_11023_n6840.n11 VSS 0.503295f
C15993 a_11023_n6840.t3 VSS 0.0377f
C15994 VDD.n0 VSS 6.14135f
C15995 VDD.n1 VSS 0.264317f
C15996 VDD.t221 VSS 0.015222f
C15997 VDD.n2 VSS 0.010908f
C15998 VDD.n3 VSS 0.010908f
C15999 VDD.n4 VSS 0.010908f
C16000 VDD.n5 VSS 0.010908f
C16001 VDD.t227 VSS 0.010959f
C16002 VDD.t220 VSS 0.071705f
C16003 VDD.t232 VSS 0.030513f
C16004 VDD.t224 VSS 0.030513f
C16005 VDD.t218 VSS 0.030513f
C16006 VDD.t230 VSS 0.030513f
C16007 VDD.t216 VSS 0.030513f
C16008 VDD.t228 VSS 0.030513f
C16009 VDD.t222 VSS 0.030513f
C16010 VDD.t234 VSS 0.030513f
C16011 VDD.t226 VSS 0.040265f
C16012 VDD.n6 VSS 0.07563f
C16013 VDD.t214 VSS 0.071705f
C16014 VDD.t206 VSS 0.030513f
C16015 VDD.t212 VSS 0.030513f
C16016 VDD.t209 VSS 0.030513f
C16017 VDD.t215 VSS 0.030513f
C16018 VDD.t211 VSS 0.030513f
C16019 VDD.t208 VSS 0.030513f
C16020 VDD.t210 VSS 0.030513f
C16021 VDD.t207 VSS 0.030513f
C16022 VDD.t213 VSS 0.040836f
C16023 VDD.n7 VSS 0.290492f
C16024 VDD.n8 VSS 0.036706f
C16025 VDD.n9 VSS 0.032972f
C16026 VDD.n10 VSS 0.032972f
C16027 VDD.n11 VSS 0.033813f
C16028 VDD.n12 VSS 0.038278f
C16029 VDD.n13 VSS 0.055661f
C16030 VDD.n14 VSS 0.100371f
C16031 VDD.t582 VSS 0.015222f
C16032 VDD.n15 VSS 0.010908f
C16033 VDD.n16 VSS 0.010908f
C16034 VDD.n17 VSS 0.010908f
C16035 VDD.n18 VSS 0.010908f
C16036 VDD.t588 VSS 0.010959f
C16037 VDD.t581 VSS 0.071705f
C16038 VDD.t593 VSS 0.030513f
C16039 VDD.t585 VSS 0.030513f
C16040 VDD.t579 VSS 0.030513f
C16041 VDD.t591 VSS 0.030513f
C16042 VDD.t577 VSS 0.030513f
C16043 VDD.t589 VSS 0.030513f
C16044 VDD.t583 VSS 0.030513f
C16045 VDD.t595 VSS 0.030513f
C16046 VDD.t587 VSS 0.040265f
C16047 VDD.n19 VSS 0.07563f
C16048 VDD.t1847 VSS 0.071705f
C16049 VDD.t1903 VSS 0.030513f
C16050 VDD.t1845 VSS 0.030513f
C16051 VDD.t1842 VSS 0.030513f
C16052 VDD.t1902 VSS 0.030513f
C16053 VDD.t1844 VSS 0.030513f
C16054 VDD.t1905 VSS 0.030513f
C16055 VDD.t1843 VSS 0.030513f
C16056 VDD.t1904 VSS 0.030513f
C16057 VDD.t1846 VSS 0.040836f
C16058 VDD.n20 VSS 0.290492f
C16059 VDD.n21 VSS 0.036706f
C16060 VDD.n22 VSS 0.032972f
C16061 VDD.n23 VSS 0.032972f
C16062 VDD.n24 VSS 0.033813f
C16063 VDD.n25 VSS 0.038278f
C16064 VDD.n26 VSS 0.079446f
C16065 VDD.t556 VSS 0.015222f
C16066 VDD.n27 VSS 0.010908f
C16067 VDD.n28 VSS 0.010908f
C16068 VDD.n29 VSS 0.010908f
C16069 VDD.n30 VSS 0.010908f
C16070 VDD.t562 VSS 0.010959f
C16071 VDD.t555 VSS 0.071705f
C16072 VDD.t567 VSS 0.030513f
C16073 VDD.t551 VSS 0.030513f
C16074 VDD.t559 VSS 0.030513f
C16075 VDD.t565 VSS 0.030513f
C16076 VDD.t553 VSS 0.030513f
C16077 VDD.t563 VSS 0.030513f
C16078 VDD.t569 VSS 0.030513f
C16079 VDD.t557 VSS 0.030513f
C16080 VDD.t561 VSS 0.040265f
C16081 VDD.n31 VSS 0.07563f
C16082 VDD.t2699 VSS 0.071705f
C16083 VDD.t2694 VSS 0.030513f
C16084 VDD.t2697 VSS 0.030513f
C16085 VDD.t2700 VSS 0.030513f
C16086 VDD.t2693 VSS 0.030513f
C16087 VDD.t2696 VSS 0.030513f
C16088 VDD.t2691 VSS 0.030513f
C16089 VDD.t2695 VSS 0.030513f
C16090 VDD.t2698 VSS 0.030513f
C16091 VDD.t2692 VSS 0.040836f
C16092 VDD.n32 VSS 0.290492f
C16093 VDD.n33 VSS 0.036706f
C16094 VDD.n34 VSS 0.032972f
C16095 VDD.n35 VSS 0.032972f
C16096 VDD.n36 VSS 0.033813f
C16097 VDD.n37 VSS 0.125281f
C16098 VDD.t668 VSS 0.015222f
C16099 VDD.n38 VSS 0.010908f
C16100 VDD.n39 VSS 0.010908f
C16101 VDD.n40 VSS 0.010908f
C16102 VDD.n41 VSS 0.010908f
C16103 VDD.t674 VSS 0.010959f
C16104 VDD.t667 VSS 0.071705f
C16105 VDD.t679 VSS 0.030513f
C16106 VDD.t683 VSS 0.030513f
C16107 VDD.t671 VSS 0.030513f
C16108 VDD.t677 VSS 0.030513f
C16109 VDD.t685 VSS 0.030513f
C16110 VDD.t675 VSS 0.030513f
C16111 VDD.t681 VSS 0.030513f
C16112 VDD.t669 VSS 0.030513f
C16113 VDD.t673 VSS 0.040265f
C16114 VDD.n42 VSS 0.07563f
C16115 VDD.t112 VSS 0.071705f
C16116 VDD.t107 VSS 0.030513f
C16117 VDD.t110 VSS 0.030513f
C16118 VDD.t113 VSS 0.030513f
C16119 VDD.t116 VSS 0.030513f
C16120 VDD.t109 VSS 0.030513f
C16121 VDD.t114 VSS 0.030513f
C16122 VDD.t108 VSS 0.030513f
C16123 VDD.t111 VSS 0.030513f
C16124 VDD.t115 VSS 0.040836f
C16125 VDD.n43 VSS 0.290492f
C16126 VDD.n44 VSS 0.036706f
C16127 VDD.n45 VSS 0.032972f
C16128 VDD.n46 VSS 0.032972f
C16129 VDD.n47 VSS 0.033813f
C16130 VDD.n48 VSS 0.042754f
C16131 VDD.n49 VSS 0.180676f
C16132 VDD.t264 VSS 0.015222f
C16133 VDD.n50 VSS 0.010908f
C16134 VDD.n51 VSS 0.010908f
C16135 VDD.n52 VSS 0.010908f
C16136 VDD.n53 VSS 0.010908f
C16137 VDD.t270 VSS 0.010959f
C16138 VDD.t263 VSS 0.071705f
C16139 VDD.t255 VSS 0.030513f
C16140 VDD.t259 VSS 0.030513f
C16141 VDD.t267 VSS 0.030513f
C16142 VDD.t253 VSS 0.030513f
C16143 VDD.t261 VSS 0.030513f
C16144 VDD.t271 VSS 0.030513f
C16145 VDD.t257 VSS 0.030513f
C16146 VDD.t265 VSS 0.030513f
C16147 VDD.t269 VSS 0.040265f
C16148 VDD.n54 VSS 0.07563f
C16149 VDD.t542 VSS 0.071705f
C16150 VDD.t547 VSS 0.030513f
C16151 VDD.t550 VSS 0.030513f
C16152 VDD.t543 VSS 0.030513f
C16153 VDD.t546 VSS 0.030513f
C16154 VDD.t549 VSS 0.030513f
C16155 VDD.t544 VSS 0.030513f
C16156 VDD.t548 VSS 0.030513f
C16157 VDD.t541 VSS 0.030513f
C16158 VDD.t545 VSS 0.040836f
C16159 VDD.n55 VSS 0.290492f
C16160 VDD.n56 VSS 0.036706f
C16161 VDD.n57 VSS 0.032972f
C16162 VDD.n58 VSS 0.032972f
C16163 VDD.n59 VSS 0.033813f
C16164 VDD.n60 VSS 0.042754f
C16165 VDD.n61 VSS 0.167887f
C16166 VDD.t1758 VSS 0.015222f
C16167 VDD.n62 VSS 0.010908f
C16168 VDD.n63 VSS 0.010908f
C16169 VDD.n64 VSS 0.010908f
C16170 VDD.n65 VSS 0.010908f
C16171 VDD.t1744 VSS 0.010959f
C16172 VDD.t1757 VSS 0.071705f
C16173 VDD.t1749 VSS 0.030513f
C16174 VDD.t1741 VSS 0.030513f
C16175 VDD.t1755 VSS 0.030513f
C16176 VDD.t1747 VSS 0.030513f
C16177 VDD.t1753 VSS 0.030513f
C16178 VDD.t1745 VSS 0.030513f
C16179 VDD.t1759 VSS 0.030513f
C16180 VDD.t1751 VSS 0.030513f
C16181 VDD.t1743 VSS 0.040265f
C16182 VDD.n66 VSS 0.07563f
C16183 VDD.t131 VSS 0.071705f
C16184 VDD.t133 VSS 0.030513f
C16185 VDD.t129 VSS 0.030513f
C16186 VDD.t136 VSS 0.030513f
C16187 VDD.t132 VSS 0.030513f
C16188 VDD.t128 VSS 0.030513f
C16189 VDD.t135 VSS 0.030513f
C16190 VDD.t127 VSS 0.030513f
C16191 VDD.t134 VSS 0.030513f
C16192 VDD.t130 VSS 0.040836f
C16193 VDD.n67 VSS 0.290492f
C16194 VDD.n68 VSS 0.036706f
C16195 VDD.n69 VSS 0.032972f
C16196 VDD.n70 VSS 0.032972f
C16197 VDD.n71 VSS 0.033813f
C16198 VDD.n72 VSS 0.042754f
C16199 VDD.n73 VSS 0.167887f
C16200 VDD.t1312 VSS 0.015222f
C16201 VDD.n74 VSS 0.010908f
C16202 VDD.n75 VSS 0.010908f
C16203 VDD.n76 VSS 0.010908f
C16204 VDD.n77 VSS 0.010908f
C16205 VDD.t1318 VSS 0.010959f
C16206 VDD.t1311 VSS 0.071705f
C16207 VDD.t1303 VSS 0.030513f
C16208 VDD.t1315 VSS 0.030513f
C16209 VDD.t1309 VSS 0.030513f
C16210 VDD.t1301 VSS 0.030513f
C16211 VDD.t1307 VSS 0.030513f
C16212 VDD.t1319 VSS 0.030513f
C16213 VDD.t1313 VSS 0.030513f
C16214 VDD.t1305 VSS 0.030513f
C16215 VDD.t1317 VSS 0.040265f
C16216 VDD.n78 VSS 0.07563f
C16217 VDD.t77 VSS 0.071705f
C16218 VDD.t79 VSS 0.030513f
C16219 VDD.t75 VSS 0.030513f
C16220 VDD.t82 VSS 0.030513f
C16221 VDD.t78 VSS 0.030513f
C16222 VDD.t74 VSS 0.030513f
C16223 VDD.t81 VSS 0.030513f
C16224 VDD.t73 VSS 0.030513f
C16225 VDD.t80 VSS 0.030513f
C16226 VDD.t76 VSS 0.040836f
C16227 VDD.n79 VSS 0.290492f
C16228 VDD.n80 VSS 0.036706f
C16229 VDD.n81 VSS 0.032972f
C16230 VDD.n82 VSS 0.032972f
C16231 VDD.n83 VSS 0.033813f
C16232 VDD.n84 VSS 0.042754f
C16233 VDD.n85 VSS 0.167887f
C16234 VDD.t98 VSS 0.015222f
C16235 VDD.n86 VSS 0.010908f
C16236 VDD.n87 VSS 0.010908f
C16237 VDD.n88 VSS 0.010908f
C16238 VDD.n89 VSS 0.010908f
C16239 VDD.t104 VSS 0.010959f
C16240 VDD.t97 VSS 0.071705f
C16241 VDD.t89 VSS 0.030513f
C16242 VDD.t101 VSS 0.030513f
C16243 VDD.t95 VSS 0.030513f
C16244 VDD.t87 VSS 0.030513f
C16245 VDD.t93 VSS 0.030513f
C16246 VDD.t105 VSS 0.030513f
C16247 VDD.t99 VSS 0.030513f
C16248 VDD.t91 VSS 0.030513f
C16249 VDD.t103 VSS 0.040265f
C16250 VDD.n90 VSS 0.07563f
C16251 VDD.t402 VSS 0.071705f
C16252 VDD.t404 VSS 0.030513f
C16253 VDD.t400 VSS 0.030513f
C16254 VDD.t407 VSS 0.030513f
C16255 VDD.t403 VSS 0.030513f
C16256 VDD.t409 VSS 0.030513f
C16257 VDD.t406 VSS 0.030513f
C16258 VDD.t408 VSS 0.030513f
C16259 VDD.t405 VSS 0.030513f
C16260 VDD.t401 VSS 0.040836f
C16261 VDD.n91 VSS 0.290492f
C16262 VDD.n92 VSS 0.036706f
C16263 VDD.n93 VSS 0.032972f
C16264 VDD.n94 VSS 0.032972f
C16265 VDD.n95 VSS 0.033813f
C16266 VDD.n96 VSS 0.042754f
C16267 VDD.n97 VSS 0.154044f
C16268 VDD.n98 VSS 0.139586f
C16269 VDD.n99 VSS 0.384295f
C16270 VDD.n100 VSS 0.047938f
C16271 VDD.n101 VSS 0.055661f
C16272 VDD.n102 VSS 0.055661f
C16273 VDD.n103 VSS 0.100371f
C16274 VDD.n104 VSS 0.100371f
C16275 VDD.n105 VSS 0.100371f
C16276 VDD.n106 VSS 0.055661f
C16277 VDD.n107 VSS 0.054895f
C16278 VDD.n108 VSS 0.346233f
C16279 VDD.n109 VSS 0.449695f
C16280 VDD.n110 VSS 0.018136f
C16281 VDD.n111 VSS 0.018136f
C16282 VDD.t373 VSS 0.02602f
C16283 VDD.n112 VSS 0.055834f
C16284 VDD.n113 VSS 0.026907f
C16285 VDD.n114 VSS 0.018136f
C16286 VDD.n115 VSS 0.018136f
C16287 VDD.t377 VSS 0.025584f
C16288 VDD.t372 VSS 0.071705f
C16289 VDD.t374 VSS 0.030513f
C16290 VDD.t378 VSS 0.030513f
C16291 VDD.t380 VSS 0.030513f
C16292 VDD.t384 VSS 0.030513f
C16293 VDD.t368 VSS 0.030513f
C16294 VDD.t382 VSS 0.030513f
C16295 VDD.t366 VSS 0.030513f
C16296 VDD.t370 VSS 0.030513f
C16297 VDD.t376 VSS 0.04154f
C16298 VDD.n116 VSS 0.096978f
C16299 VDD.n117 VSS 0.030194f
C16300 VDD.n118 VSS 0.023996f
C16301 VDD.n119 VSS 0.053197f
C16302 VDD.n120 VSS 0.275749f
C16303 VDD.n122 VSS 0.073678f
C16304 VDD.n124 VSS 0.380204f
C16305 VDD.n126 VSS 0.073678f
C16306 VDD.n128 VSS 0.055258f
C16307 VDD.n129 VSS 0.268995f
C16308 VDD.t843 VSS 0.083207f
C16309 VDD.n130 VSS 0.01095f
C16310 VDD.n131 VSS 0.268995f
C16311 VDD.t2021 VSS 0.081486f
C16312 VDD.t2022 VSS 0.012817f
C16313 VDD.n132 VSS 0.065636f
C16314 VDD.t2351 VSS 0.081486f
C16315 VDD.t2352 VSS 0.012812f
C16316 VDD.n133 VSS 0.066773f
C16317 VDD.n134 VSS 0.021593f
C16318 VDD.n135 VSS 0.016238f
C16319 VDD.n136 VSS 0.268995f
C16320 VDD.n137 VSS 0.01095f
C16321 VDD.n138 VSS 0.268995f
C16322 VDD.t436 VSS 0.083544f
C16323 VDD.n139 VSS 0.083549f
C16324 VDD.n140 VSS 0.268995f
C16325 VDD.n141 VSS 0.01095f
C16326 VDD.t2009 VSS 0.081468f
C16327 VDD.t2010 VSS 0.011814f
C16328 VDD.n142 VSS 0.076553f
C16329 VDD.t2011 VSS 0.081468f
C16330 VDD.t2012 VSS 0.011792f
C16331 VDD.n143 VSS 0.073782f
C16332 VDD.n144 VSS 0.025123f
C16333 VDD.n145 VSS 0.029497f
C16334 VDD.n146 VSS 0.01095f
C16335 VDD.n147 VSS 0.268995f
C16336 VDD.n148 VSS 0.268995f
C16337 VDD.n149 VSS 0.268995f
C16338 VDD.n150 VSS 0.01095f
C16339 VDD.n151 VSS 0.01095f
C16340 VDD.n153 VSS 0.268995f
C16341 VDD.n154 VSS 0.268995f
C16342 VDD.n156 VSS 0.01095f
C16343 VDD.n157 VSS 0.01095f
C16344 VDD.n158 VSS 0.268995f
C16345 VDD.n159 VSS 0.268995f
C16346 VDD.n160 VSS 0.268995f
C16347 VDD.n161 VSS 0.01095f
C16348 VDD.n162 VSS 0.01095f
C16349 VDD.n164 VSS 0.268995f
C16350 VDD.n165 VSS 0.268995f
C16351 VDD.n167 VSS 0.01095f
C16352 VDD.n168 VSS 0.01095f
C16353 VDD.n169 VSS 0.268995f
C16354 VDD.n170 VSS 0.268995f
C16355 VDD.n171 VSS 0.268995f
C16356 VDD.n172 VSS 0.01095f
C16357 VDD.n173 VSS 0.01095f
C16358 VDD.n174 VSS 0.0761f
C16359 VDD.n175 VSS 0.711807f
C16360 VDD.n176 VSS 0.016025f
C16361 VDD.n177 VSS 0.016025f
C16362 VDD.t340 VSS 0.023024f
C16363 VDD.t331 VSS 0.071705f
C16364 VDD.t329 VSS 0.030513f
C16365 VDD.t333 VSS 0.030513f
C16366 VDD.t327 VSS 0.030513f
C16367 VDD.t325 VSS 0.030513f
C16368 VDD.t345 VSS 0.030513f
C16369 VDD.t343 VSS 0.030513f
C16370 VDD.t337 VSS 0.030513f
C16371 VDD.t341 VSS 0.030513f
C16372 VDD.t339 VSS 0.041137f
C16373 VDD.n178 VSS 0.091674f
C16374 VDD.n179 VSS 0.028342f
C16375 VDD.n180 VSS 0.021061f
C16376 VDD.n181 VSS 0.016025f
C16377 VDD.n182 VSS 0.016025f
C16378 VDD.t332 VSS 0.023567f
C16379 VDD.n183 VSS 0.050956f
C16380 VDD.n184 VSS 0.025638f
C16381 VDD.n186 VSS 0.232747f
C16382 VDD.n187 VSS 0.686399f
C16383 VDD.n188 VSS -0.054026f
C16384 VDD.n190 VSS 0.073678f
C16385 VDD.n191 VSS 0.073678f
C16386 VDD.n192 VSS 0.073678f
C16387 VDD.n196 VSS 0.073678f
C16388 VDD.n197 VSS 0.073678f
C16389 VDD.n198 VSS 0.380204f
C16390 VDD.n199 VSS 0.044796f
C16391 VDD.n200 VSS 0.044796f
C16392 VDD.n202 VSS 0.073678f
C16393 VDD.n203 VSS 0.073678f
C16394 VDD.n204 VSS 0.073678f
C16395 VDD.n208 VSS 0.073678f
C16396 VDD.n209 VSS 0.073678f
C16397 VDD.n210 VSS 0.055258f
C16398 VDD.n211 VSS -0.055518f
C16399 VDD.n212 VSS 5.12404f
C16400 VDD.n213 VSS 21.3749f
C16401 VDD.n214 VSS 0.302928f
C16402 VDD.n215 VSS 0.429013f
C16403 VDD.n216 VSS 0.118404f
C16404 VDD.t2048 VSS 0.07726f
C16405 VDD.t1162 VSS 0.088298f
C16406 VDD.t2792 VSS 0.088298f
C16407 VDD.t2218 VSS 0.088298f
C16408 VDD.t2086 VSS 0.088298f
C16409 VDD.t1461 VSS 0.088298f
C16410 VDD.t1002 VSS 0.088298f
C16411 VDD.t2094 VSS 0.07726f
C16412 VDD.n218 VSS 0.04743f
C16413 VDD.t2236 VSS 0.033112f
C16414 VDD.t2046 VSS 0.033112f
C16415 VDD.n219 VSS 0.04743f
C16416 VDD.n220 VSS 0.015305f
C16417 VDD.n221 VSS 0.118404f
C16418 VDD.t2811 VSS 0.069504f
C16419 VDD.t2894 VSS 0.044149f
C16420 VDD.t3830 VSS 0.044149f
C16421 VDD.t3827 VSS 0.044149f
C16422 VDD.t3305 VSS 0.044149f
C16423 VDD.t1945 VSS 0.044149f
C16424 VDD.t904 VSS 0.044149f
C16425 VDD.t1634 VSS 0.044149f
C16426 VDD.t3778 VSS 0.044149f
C16427 VDD.t3166 VSS 0.044149f
C16428 VDD.t3877 VSS 0.044149f
C16429 VDD.t1898 VSS 0.044149f
C16430 VDD.t874 VSS 0.044149f
C16431 VDD.t1280 VSS 0.044149f
C16432 VDD.t3171 VSS 0.044149f
C16433 VDD.t1103 VSS 0.044149f
C16434 VDD.t2516 VSS 0.044149f
C16435 VDD.t3943 VSS 0.069504f
C16436 VDD.t2468 VSS 0.044149f
C16437 VDD.t2271 VSS 0.044149f
C16438 VDD.t1105 VSS 0.044149f
C16439 VDD.t2203 VSS 0.044149f
C16440 VDD.t3314 VSS 0.044149f
C16441 VDD.t2153 VSS 0.044149f
C16442 VDD.t3180 VSS 0.044149f
C16443 VDD.t2090 VSS 0.044149f
C16444 VDD.t1575 VSS 0.044149f
C16445 VDD.t2220 VSS 0.044149f
C16446 VDD.t2472 VSS 0.044149f
C16447 VDD.t2273 VSS 0.044149f
C16448 VDD.t3169 VSS 0.044149f
C16449 VDD.t2264 VSS 0.044149f
C16450 VDD.t3146 VSS 0.044149f
C16451 VDD.t2571 VSS 0.044149f
C16452 VDD.t2510 VSS 0.080541f
C16453 VDD.t2455 VSS 0.066223f
C16454 VDD.t2796 VSS 0.044149f
C16455 VDD.t2837 VSS 0.044149f
C16456 VDD.t2487 VSS 0.044149f
C16457 VDD.t4236 VSS 0.044149f
C16458 VDD.t2115 VSS 0.044149f
C16459 VDD.t3301 VSS 0.044149f
C16460 VDD.t3875 VSS 0.044149f
C16461 VDD.t1441 VSS 0.02917f
C16462 VDD.t4062 VSS 0.044149f
C16463 VDD.t2457 VSS 0.070165f
C16464 VDD.t1142 VSS 0.044149f
C16465 VDD.t1988 VSS 0.044149f
C16466 VDD.t2174 VSS 0.044149f
C16467 VDD.t1969 VSS 0.044149f
C16468 VDD.t3538 VSS 0.080541f
C16469 VDD.t1584 VSS 0.088298f
C16470 VDD.t1607 VSS 0.088298f
C16471 VDD.t3554 VSS 0.088298f
C16472 VDD.t3335 VSS 0.088298f
C16473 VDD.t3343 VSS 0.088298f
C16474 VDD.t1239 VSS 0.088298f
C16475 VDD.t1609 VSS 0.088298f
C16476 VDD.t908 VSS 0.078178f
C16477 VDD.n223 VSS 0.121999f
C16478 VDD.n224 VSS 0.019165f
C16479 VDD.n225 VSS 0.019165f
C16480 VDD.n226 VSS 0.019165f
C16481 VDD.n227 VSS 0.019165f
C16482 VDD.n228 VSS 0.019165f
C16483 VDD.n229 VSS 0.014594f
C16484 VDD.n230 VSS 0.118404f
C16485 VDD.n231 VSS 0.014557f
C16486 VDD.t2599 VSS 0.047105f
C16487 VDD.t2099 VSS 0.035674f
C16488 VDD.t4111 VSS 0.036955f
C16489 VDD.t2544 VSS 0.044149f
C16490 VDD.t205 VSS 0.020103f
C16491 VDD.t4112 VSS 0.043163f
C16492 VDD.t349 VSS 0.043262f
C16493 VDD.t472 VSS 0.036364f
C16494 VDD.t634 VSS 0.055186f
C16495 VDD.t4122 VSS 0.020103f
C16496 VDD.t4057 VSS 0.044149f
C16497 VDD.t641 VSS 0.044839f
C16498 VDD.t2464 VSS 0.02917f
C16499 VDD.t3200 VSS 0.046317f
C16500 VDD.t777 VSS 0.044149f
C16501 VDD.t3269 VSS 0.037053f
C16502 VDD.t1769 VSS 0.040207f
C16503 VDD.t642 VSS 0.033112f
C16504 VDD.t1054 VSS 0.026016f
C16505 VDD.n238 VSS 0.04743f
C16506 VDD.n240 VSS 0.118404f
C16507 VDD.n243 VSS 0.012831f
C16508 VDD.t3144 VSS 0.07726f
C16509 VDD.t2385 VSS 0.088298f
C16510 VDD.t1328 VSS 0.088298f
C16511 VDD.t1201 VSS 0.088298f
C16512 VDD.t953 VSS 0.088298f
C16513 VDD.t2366 VSS 0.088298f
C16514 VDD.t2776 VSS 0.088298f
C16515 VDD.t988 VSS 0.088298f
C16516 VDD.t3644 VSS 0.080541f
C16517 VDD.n252 VSS 0.118404f
C16518 VDD.t3626 VSS 0.080541f
C16519 VDD.t2323 VSS 0.088298f
C16520 VDD.t2266 VSS 0.088298f
C16521 VDD.t2147 VSS 0.088298f
C16522 VDD.t1368 VSS 0.088298f
C16523 VDD.t1419 VSS 0.081202f
C16524 VDD.t496 VSS 0.044149f
C16525 VDD.t4139 VSS 0.048288f
C16526 VDD.t281 VSS 0.044149f
C16527 VDD.t4078 VSS 0.020103f
C16528 VDD.t1726 VSS 0.044149f
C16529 VDD.t2727 VSS 0.034294f
C16530 VDD.t1413 VSS 0.027396f
C16531 VDD.t3991 VSS 0.025819f
C16532 VDD.n255 VSS 0.023384f
C16533 VDD.t1729 VSS 0.033604f
C16534 VDD.t3127 VSS 0.020103f
C16535 VDD.t3526 VSS 0.022074f
C16536 VDD.t1578 VSS 0.031141f
C16537 VDD.t534 VSS 0.016556f
C16538 VDD.t1577 VSS 0.034382f
C16539 VDD.t2078 VSS 0.043682f
C16540 VDD.t2480 VSS 0.027876f
C16541 VDD.t1728 VSS 0.016038f
C16542 VDD.t2478 VSS 0.0287f
C16543 VDD.t3990 VSS 0.032475f
C16544 VDD.t3612 VSS 0.020103f
C16545 VDD.t1624 VSS 0.036659f
C16546 VDD.t511 VSS 0.035181f
C16547 VDD.t466 VSS 0.020103f
C16548 VDD.t2503 VSS 0.043656f
C16549 VDD.t1622 VSS 0.034787f
C16550 VDD.t530 VSS 0.037053f
C16551 VDD.t3650 VSS 0.047795f
C16552 VDD.t2685 VSS 0.020103f
C16553 VDD.t3150 VSS 0.028973f
C16554 VDD.t3597 VSS 0.025425f
C16555 VDD.t2564 VSS 0.020103f
C16556 VDD.t1837 VSS 0.020103f
C16557 VDD.t525 VSS 0.029761f
C16558 VDD.t2683 VSS 0.026312f
C16559 VDD.n262 VSS 0.023385f
C16560 VDD.t3919 VSS 0.030225f
C16561 VDD.t2258 VSS 0.029651f
C16562 VDD.t1959 VSS 0.019475f
C16563 VDD.t775 VSS 0.022435f
C16564 VDD.t631 VSS 0.024917f
C16565 VDD.t1977 VSS 0.035449f
C16566 VDD.t2231 VSS 0.034405f
C16567 VDD.t490 VSS 0.03252f
C16568 VDD.t2459 VSS 0.031141f
C16569 VDD.t1356 VSS 0.016556f
C16570 VDD.t2461 VSS 0.020103f
C16571 VDD.t1962 VSS 0.025819f
C16572 VDD.t3920 VSS 0.037251f
C16573 VDD.t1211 VSS 0.020103f
C16574 VDD.t2466 VSS 0.016556f
C16575 VDD.t1209 VSS 0.034294f
C16576 VDD.t1960 VSS 0.027987f
C16577 VDD.t4258 VSS 0.020103f
C16578 VDD.t2624 VSS 0.016556f
C16579 VDD.t4257 VSS 0.044149f
C16580 VDD.t3275 VSS 0.042966f
C16581 VDD.t1183 VSS 0.019118f
C16582 VDD.t1184 VSS 0.021483f
C16583 VDD.t3487 VSS 0.022074f
C16584 VDD.t1140 VSS 0.020103f
C16585 VDD.t2968 VSS 0.044149f
C16586 VDD.n269 VSS 0.063099f
C16587 VDD.t1571 VSS 0.045528f
C16588 VDD.t3980 VSS 0.034294f
C16589 VDD.t4216 VSS 0.023651f
C16590 VDD.t1261 VSS 0.020103f
C16591 VDD.t469 VSS 0.028283f
C16592 VDD.t1569 VSS 0.032422f
C16593 VDD.t3741 VSS 0.020103f
C16594 VDD.t3849 VSS 0.022074f
C16595 VDD.t3743 VSS 0.029602f
C16596 VDD.t2140 VSS 0.020896f
C16597 VDD.t3737 VSS 0.023676f
C16598 VDD.t3739 VSS 0.025585f
C16599 VDD.t3791 VSS 0.021353f
C16600 VDD.t1875 VSS 0.034252f
C16601 VDD.t497 VSS 0.022074f
C16602 VDD.t1920 VSS 0.027593f
C16603 VDD.t2003 VSS 0.025622f
C16604 VDD.t3850 VSS 0.022074f
C16605 VDD.t2001 VSS 0.020103f
C16606 VDD.t2141 VSS 0.02168f
C16607 VDD.t3848 VSS 0.020498f
C16608 VDD.t1918 VSS 0.020103f
C16609 VDD.t1533 VSS 0.022074f
C16610 VDD.t1877 VSS 0.02444f
C16611 VDD.t1873 VSS 0.031929f
C16612 VDD.t2138 VSS 0.022074f
C16613 VDD.t2005 VSS 0.020103f
C16614 VDD.t2628 VSS 0.038942f
C16615 VDD.n279 VSS 0.105436f
C16616 VDD.n283 VSS 0.012965f
C16617 VDD.n288 VSS 0.013184f
C16618 VDD.n289 VSS 0.010869f
C16619 VDD.n291 VSS 0.118404f
C16620 VDD.t3692 VSS 0.031633f
C16621 VDD.t1838 VSS 0.037251f
C16622 VDD.t2543 VSS 0.024932f
C16623 VDD.t3600 VSS 0.020103f
C16624 VDD.t3106 VSS 0.023651f
C16625 VDD.t2076 VSS 0.020103f
C16626 VDD.t3212 VSS 0.041685f
C16627 VDD.t4240 VSS 0.037053f
C16628 VDD.t2057 VSS 0.022074f
C16629 VDD.t3175 VSS 0.031535f
C16630 VDD.t3177 VSS 0.019315f
C16631 VDD.t3887 VSS 0.022863f
C16632 VDD.t494 VSS 0.042178f
C16633 VDD.t2853 VSS 0.02444f
C16634 VDD.t2059 VSS 0.016556f
C16635 VDD.t2854 VSS 0.020103f
C16636 VDD.t2082 VSS 0.032436f
C16637 VDD.t2550 VSS 0.028678f
C16638 VDD.t1504 VSS 0.030836f
C16639 VDD.t2989 VSS 0.045995f
C16640 VDD.t465 VSS 0.034271f
C16641 VDD.t483 VSS 0.046711f
C16642 VDD.t3772 VSS 0.039616f
C16643 VDD.t323 VSS 0.020103f
C16644 VDD.t1505 VSS 0.026016f
C16645 VDD.n303 VSS 0.023385f
C16646 VDD.n308 VSS 0.118404f
C16647 VDD.t4179 VSS 0.029257f
C16648 VDD.t3089 VSS 0.026731f
C16649 VDD.t1497 VSS 0.020621f
C16650 VDD.t1278 VSS 0.021845f
C16651 VDD.t2847 VSS 0.030661f
C16652 VDD.t3749 VSS 0.026903f
C16653 VDD.t1519 VSS 0.044247f
C16654 VDD.t4059 VSS 0.02444f
C16655 VDD.t729 VSS 0.020399f
C16656 VDD.t3466 VSS 0.022764f
C16657 VDD.t4154 VSS 0.034294f
C16658 VDD.t1517 VSS 0.040601f
C16659 VDD.t3499 VSS 0.032619f
C16660 VDD.t1465 VSS 0.032323f
C16661 VDD.t2474 VSS 0.033112f
C16662 VDD.t4152 VSS 0.039616f
C16663 VDD.t731 VSS 0.036955f
C16664 VDD.t895 VSS 0.041882f
C16665 VDD.t9 VSS 0.02237f
C16666 VDD.t522 VSS 0.03932f
C16667 VDD.t1132 VSS 0.044149f
C16668 VDD.t3 VSS 0.044149f
C16669 VDD.t3204 VSS 0.073446f
C16670 VDD.n319 VSS 0.118404f
C16671 VDD.t2370 VSS 0.073446f
C16672 VDD.t4117 VSS 0.044149f
C16673 VDD.t2753 VSS 0.044149f
C16674 VDD.t4060 VSS 0.03932f
C16675 VDD.t4109 VSS 0.02237f
C16676 VDD.t1771 VSS 0.041882f
C16677 VDD.t639 VSS 0.035083f
C16678 VDD.t1066 VSS 0.033407f
C16679 VDD.t3858 VSS 0.041882f
C16680 VDD.t4061 VSS 0.034984f
C16681 VDD.t649 VSS 0.02306f
C16682 VDD.t413 VSS 0.02306f
C16683 VDD.t3985 VSS 0.036265f
C16684 VDD.t1796 VSS 0.046711f
C16685 VDD.t1475 VSS 0.055186f
C16686 VDD.t1774 VSS 0.040601f
C16687 VDD.t790 VSS 0.023651f
C16688 VDD.t1871 VSS 0.025819f
C16689 VDD.t1050 VSS 0.033309f
C16690 VDD.t1052 VSS 0.033604f
C16691 VDD.t1118 VSS 0.034294f
C16692 VDD.n325 VSS 0.035801f
C16693 VDD.t3517 VSS 0.026312f
C16694 VDD.t3519 VSS 0.045923f
C16695 VDD.t2841 VSS 0.044937f
C16696 VDD.t2144 VSS 0.022074f
C16697 VDD.t2655 VSS 0.016556f
C16698 VDD.t2145 VSS 0.016556f
C16699 VDD.t2654 VSS 0.022074f
C16700 VDD.t2040 VSS 0.044937f
C16701 VDD.t2211 VSS 0.045923f
C16702 VDD.t2212 VSS 0.027494f
C16703 VDD.t3675 VSS 0.03252f
C16704 VDD.t3955 VSS 0.022074f
C16705 VDD.t3677 VSS 0.026312f
C16706 VDD.t2530 VSS 0.051047f
C16707 VDD.t2595 VSS 0.034688f
C16708 VDD.t646 VSS 0.023651f
C16709 VDD.t4284 VSS 0.020103f
C16710 VDD.t3825 VSS 0.026016f
C16711 VDD.t3864 VSS 0.036659f
C16712 VDD.t4209 VSS 0.020103f
C16713 VDD.t3860 VSS 0.023651f
C16714 VDD.t1056 VSS 0.040207f
C16715 VDD.t651 VSS 0.052821f
C16716 VDD.t1916 VSS 0.036462f
C16717 VDD.n334 VSS 0.023385f
C16718 VDD.n342 VSS 0.126498f
C16719 VDD.t1022 VSS 0.253425f
C16720 VDD.t2279 VSS 0.011964f
C16721 VDD.t513 VSS 0.02556f
C16722 VDD.t2926 VSS 0.034805f
C16723 VDD.t955 VSS 0.061997f
C16724 VDD.t238 VSS 0.032514f
C16725 VDD.t1795 VSS 0.026764f
C16726 VDD.n348 VSS 0.079196f
C16727 VDD.t2374 VSS 0.092286f
C16728 VDD.t786 VSS 0.027901f
C16729 VDD.t1930 VSS 0.037524f
C16730 VDD.n349 VSS 0.012601f
C16731 VDD.t996 VSS 0.05112f
C16732 VDD.n350 VSS 0.068049f
C16733 VDD.t1931 VSS 0.018043f
C16734 VDD.t3951 VSS 0.031504f
C16735 VDD.t4070 VSS 0.027876f
C16736 VDD.t3669 VSS 0.02757f
C16737 VDD.t533 VSS 0.034271f
C16738 VDD.t473 VSS 0.046711f
C16739 VDD.t3182 VSS 0.036462f
C16740 VDD.t1267 VSS 0.020103f
C16741 VDD.t3954 VSS 0.034885f
C16742 VDD.t3785 VSS 0.040207f
C16743 VDD.t2922 VSS 0.02444f
C16744 VDD.t1095 VSS 0.02444f
C16745 VDD.t3489 VSS 0.029958f
C16746 VDD.t3952 VSS 0.024045f
C16747 VDD.t2740 VSS 0.020103f
C16748 VDD.t2632 VSS 0.036967f
C16749 VDD.n351 VSS 0.104042f
C16750 VDD.n353 VSS 0.010131f
C16751 VDD.n354 VSS 0.014137f
C16752 VDD.n355 VSS 0.017063f
C16753 VDD.n356 VSS 0.013846f
C16754 VDD.n357 VSS 0.015669f
C16755 VDD.n358 VSS 0.012481f
C16756 VDD.n359 VSS 0.118404f
C16757 VDD.t3192 VSS 0.040207f
C16758 VDD.t506 VSS 0.063267f
C16759 VDD.t4046 VSS 0.055186f
C16760 VDD.t4120 VSS 0.022074f
C16761 VDD.t1114 VSS 0.032028f
C16762 VDD.t1113 VSS 0.020892f
C16763 VDD.t2928 VSS 0.036856f
C16764 VDD.t980 VSS 0.040601f
C16765 VDD.t2454 VSS 0.016556f
C16766 VDD.t979 VSS 0.016556f
C16767 VDD.t2452 VSS 0.040601f
C16768 VDD.t2886 VSS 0.036856f
C16769 VDD.t2879 VSS 0.020892f
C16770 VDD.t2880 VSS 0.03863f
C16771 VDD.t1326 VSS 0.029663f
C16772 VDD.t633 VSS 0.049569f
C16773 VDD.t1082 VSS 0.077457f
C16774 VDD.t3580 VSS 0.046317f
C16775 VDD.t637 VSS 0.020103f
C16776 VDD.t440 VSS 0.02695f
C16777 VDD.n373 VSS 0.031182f
C16778 VDD.n379 VSS 0.118404f
C16779 VDD.n381 VSS 0.010563f
C16780 VDD.t611 VSS 0.034491f
C16781 VDD.t173 VSS 0.045331f
C16782 VDD.t149 VSS 0.022074f
C16783 VDD.t171 VSS 0.024045f
C16784 VDD.t145 VSS 0.022074f
C16785 VDD.t175 VSS 0.020103f
C16786 VDD.t153 VSS 0.022074f
C16787 VDD.t177 VSS 0.024045f
C16788 VDD.t147 VSS 0.022074f
C16789 VDD.t187 VSS 0.023651f
C16790 VDD.t841 VSS 0.022074f
C16791 VDD.t161 VSS 0.024045f
C16792 VDD.t831 VSS 0.022074f
C16793 VDD.t157 VSS 0.020103f
C16794 VDD.t837 VSS 0.022074f
C16795 VDD.t159 VSS 0.024045f
C16796 VDD.t833 VSS 0.022074f
C16797 VDD.t167 VSS 0.020103f
C16798 VDD.t827 VSS 0.022074f
C16799 VDD.t163 VSS 0.024045f
C16800 VDD.t839 VSS 0.022074f
C16801 VDD.t169 VSS 0.020103f
C16802 VDD.t829 VSS 0.022074f
C16803 VDD.t165 VSS 0.024045f
C16804 VDD.t835 VSS 0.022074f
C16805 VDD.t179 VSS 0.022863f
C16806 VDD.t183 VSS 0.03794f
C16807 VDD.t1036 VSS 0.022074f
C16808 VDD.t181 VSS 0.020103f
C16809 VDD.t3094 VSS 0.022074f
C16810 VDD.t185 VSS 0.028874f
C16811 VDD.n401 VSS 0.028903f
C16812 VDD.n406 VSS 0.118404f
C16813 VDD.n407 VSS 0.011854f
C16814 VDD.n409 VSS 0.023385f
C16815 VDD.t4092 VSS 0.030155f
C16816 VDD.t335 VSS 0.024045f
C16817 VDD.t4086 VSS 0.023651f
C16818 VDD.t3228 VSS 0.020103f
C16819 VDD.t4090 VSS 0.024834f
C16820 VDD.t4094 VSS 0.041784f
C16821 VDD.t1166 VSS 0.023651f
C16822 VDD.t821 VSS 0.023651f
C16823 VDD.t2882 VSS 0.024045f
C16824 VDD.t817 VSS 0.02641f
C16825 VDD.t819 VSS 0.036265f
C16826 VDD.t4127 VSS 0.024045f
C16827 VDD.t825 VSS 0.020103f
C16828 VDD.t3551 VSS 0.034294f
C16829 VDD.t3698 VSS 0.034294f
C16830 VDD.t39 VSS 0.032323f
C16831 VDD.t2813 VSS 0.040207f
C16832 VDD.t1079 VSS 0.040207f
C16833 VDD.t35 VSS 0.040207f
C16834 VDD.t3390 VSS 0.031141f
C16835 VDD.t701 VSS 0.020103f
C16836 VDD.t3394 VSS 0.02925f
C16837 VDD.t30 VSS 0.024679f
C16838 VDD.t2964 VSS 0.019475f
C16839 VDD.t3735 VSS 0.027876f
C16840 VDD.t3553 VSS 0.027685f
C16841 VDD.n420 VSS 0.032182f
C16842 VDD.t2814 VSS 0.035043f
C16843 VDD.t1527 VSS 0.033801f
C16844 VDD.t2723 VSS 0.02444f
C16845 VDD.t706 VSS 0.02444f
C16846 VDD.t1168 VSS 0.020103f
C16847 VDD.t2524 VSS 0.020103f
C16848 VDD.t2978 VSS 0.034294f
C16849 VDD.t1529 VSS 0.034294f
C16850 VDD.t24 VSS 0.020103f
C16851 VDD.t1531 VSS 0.020103f
C16852 VDD.t1048 VSS 0.043251f
C16853 VDD.t1040 VSS 0.031514f
C16854 VDD.t4026 VSS 0.019522f
C16855 VDD.t37 VSS 0.034067f
C16856 VDD.t32 VSS 0.020287f
C16857 VDD.t2054 VSS 0.019522f
C16858 VDD.t1038 VSS 0.019522f
C16859 VDD.t1084 VSS 0.020287f
C16860 VDD.t617 VSS 0.026389f
C16861 VDD.t1042 VSS 0.020869f
C16862 VDD.t807 VSS 0.020103f
C16863 VDD.t26 VSS 0.020103f
C16864 VDD.t813 VSS 0.020103f
C16865 VDD.t1086 VSS 0.020103f
C16866 VDD.t597 VSS 0.020103f
C16867 VDD.t1060 VSS 0.020103f
C16868 VDD.t1088 VSS 0.020103f
C16869 VDD.t1058 VSS 0.020103f
C16870 VDD.t2050 VSS 0.020103f
C16871 VDD.t1090 VSS 0.027987f
C16872 VDD.t1075 VSS 0.020301f
C16873 VDD.n432 VSS 0.023385f
C16874 VDD.t1062 VSS 0.031633f
C16875 VDD.t1870 VSS 0.020103f
C16876 VDD.t3823 VSS 0.020103f
C16877 VDD.t3757 VSS 0.020103f
C16878 VDD.t3731 VSS 0.020103f
C16879 VDD.t3817 VSS 0.03183f
C16880 VDD.t3021 VSS 0.046612f
C16881 VDD.t3844 VSS 0.041882f
C16882 VDD.t2180 VSS 0.03252f
C16883 VDD.t1155 VSS 0.023651f
C16884 VDD.t3244 VSS 0.016556f
C16885 VDD.t1157 VSS 0.053018f
C16886 VDD.t1398 VSS 0.059522f
C16887 VDD.t1399 VSS 0.020596f
C16888 VDD.t2851 VSS 0.027987f
C16889 VDD.t1885 VSS 0.03252f
C16890 VDD.t2593 VSS 0.016556f
C16891 VDD.t1884 VSS 0.016556f
C16892 VDD.t2592 VSS 0.042966f
C16893 VDD.t3760 VSS 0.044937f
C16894 VDD.t1336 VSS 0.016556f
C16895 VDD.t3761 VSS 0.016556f
C16896 VDD.t1334 VSS 0.022074f
C16897 VDD.t3758 VSS 0.022074f
C16898 VDD.t2246 VSS 0.033112f
C16899 VDD.n441 VSS 0.044473f
C16900 VDD.t1859 VSS 0.038039f
C16901 VDD.t1892 VSS 0.034294f
C16902 VDD.t2015 VSS 0.020103f
C16903 VDD.t1325 VSS 0.020103f
C16904 VDD.t463 VSS 0.022074f
C16905 VDD.t3498 VSS 0.02444f
C16906 VDD.t1861 VSS 0.022074f
C16907 VDD.t1064 VSS 0.020103f
C16908 VDD.t3264 VSS 0.037543f
C16909 VDD.t925 VSS 0.028732f
C16910 VDD.t1715 VSS 0.019475f
C16911 VDD.t3104 VSS 0.027876f
C16912 VDD.t2970 VSS 0.019475f
C16913 VDD.t2240 VSS 0.023564f
C16914 VDD.t1266 VSS 0.030331f
C16915 VDD.t527 VSS 0.039714f
C16916 VDD.t4141 VSS 0.031141f
C16917 VDD.t3331 VSS 0.020103f
C16918 VDD.t3488 VSS 0.020103f
C16919 VDD.t1714 VSS 0.02168f
C16920 VDD.t3265 VSS 0.022469f
C16921 VDD.t2518 VSS 0.020103f
C16922 VDD.t1027 VSS 0.048485f
C16923 VDD.t2065 VSS 0.034294f
C16924 VDD.t1716 VSS 0.023651f
C16925 VDD.t398 VSS 0.051188f
C16926 VDD.n447 VSS 0.112724f
C16927 VDD.n448 VSS 0.010268f
C16928 VDD.n449 VSS 0.0137f
C16929 VDD.n450 VSS 0.011673f
C16930 VDD.n452 VSS 0.012997f
C16931 VDD.n453 VSS 0.011158f
C16932 VDD.n454 VSS 0.01306f
C16933 VDD.n456 VSS 0.118404f
C16934 VDD.t3892 VSS 0.044881f
C16935 VDD.t2355 VSS 0.028709f
C16936 VDD.t1164 VSS 0.030622f
C16937 VDD.t3482 VSS 0.037512f
C16938 VDD.t3481 VSS 0.017225f
C16939 VDD.t504 VSS 0.020636f
C16940 VDD.t4230 VSS 0.043709f
C16941 VDD.t1613 VSS 0.031141f
C16942 VDD.t3632 VSS 0.016556f
C16943 VDD.t1614 VSS 0.017738f
C16944 VDD.t2358 VSS 0.03252f
C16945 VDD.t4234 VSS 0.024932f
C16946 VDD.t3891 VSS 0.021188f
C16947 VDD.t3327 VSS 0.043755f
C16948 VDD.t1282 VSS 0.038236f
C16949 VDD.t2356 VSS 0.023651f
C16950 VDD.t3776 VSS 0.020103f
C16951 VDD.t394 VSS 0.053412f
C16952 VDD.t3256 VSS 0.061789f
C16953 VDD.t4114 VSS 0.022074f
C16954 VDD.t3254 VSS 0.020103f
C16955 VDD.t1230 VSS 0.025819f
C16956 VDD.t3720 VSS 0.020103f
C16957 VDD.t3925 VSS 0.028184f
C16958 VDD.n473 VSS 0.023385f
C16959 VDD.n480 VSS 0.118404f
C16960 VDD.n482 VSS 0.010149f
C16961 VDD.t7 VSS 0.033604f
C16962 VDD.t605 VSS 0.025819f
C16963 VDD.t1274 VSS 0.022074f
C16964 VDD.t1954 VSS 0.022074f
C16965 VDD.t1272 VSS 0.016556f
C16966 VDD.t1953 VSS 0.052131f
C16967 VDD.t3443 VSS 0.049667f
C16968 VDD.t2541 VSS 0.016556f
C16969 VDD.t3444 VSS 0.022074f
C16970 VDD.t1347 VSS 0.026805f
C16971 VDD.t1349 VSS 0.022271f
C16972 VDD.t2319 VSS 0.044937f
C16973 VDD.t1395 VSS 0.044839f
C16974 VDD.t3121 VSS 0.016556f
C16975 VDD.t1396 VSS 0.023651f
C16976 VDD.t3606 VSS 0.03252f
C16977 VDD.t2862 VSS 0.049273f
C16978 VDD.t1508 VSS 0.050554f
C16979 VDD.t725 VSS 0.023651f
C16980 VDD.t3026 VSS 0.044149f
C16981 VDD.t519 VSS 0.046908f
C16982 VDD.t2805 VSS 0.027396f
C16983 VDD.t2803 VSS 0.031732f
C16984 VDD.n494 VSS 0.028903f
C16985 VDD.n499 VSS 0.231769f
C16986 VDD.n502 VSS 0.029197f
C16987 VDD.t732 VSS 0.033785f
C16988 VDD.t747 VSS 0.038827f
C16989 VDD.t2784 VSS 0.047499f
C16990 VDD.t717 VSS 0.020103f
C16991 VDD.t2986 VSS 0.023848f
C16992 VDD.t4013 VSS 0.040207f
C16993 VDD.t3307 VSS 0.026706f
C16994 VDD.t418 VSS 0.034294f
C16995 VDD.t2984 VSS 0.03252f
C16996 VDD.t2104 VSS 0.020103f
C16997 VDD.t4129 VSS 0.016556f
C16998 VDD.t2103 VSS 0.037251f
C16999 VDD.t1853 VSS 0.044937f
C17000 VDD.t3446 VSS 0.021089f
C17001 VDD.t1855 VSS 0.016556f
C17002 VDD.t3447 VSS 0.024045f
C17003 VDD.t2976 VSS 0.022074f
C17004 VDD.t1544 VSS 0.025228f
C17005 VDD.t4262 VSS 0.042868f
C17006 VDD.t3033 VSS 0.02237f
C17007 VDD.t2186 VSS 0.014585f
C17008 VDD.t3801 VSS 0.022074f
C17009 VDD.t3054 VSS 0.020103f
C17010 VDD.t3031 VSS 0.016556f
C17011 VDD.t3053 VSS 0.044346f
C17012 VDD.n510 VSS 0.048218f
C17013 VDD.t4250 VSS 0.023355f
C17014 VDD.t4251 VSS 0.032422f
C17015 VDD.t20 VSS 0.03252f
C17016 VDD.t1767 VSS 0.025819f
C17017 VDD.t1392 VSS 0.031239f
C17018 VDD.t1390 VSS 0.027199f
C17019 VDD.t743 VSS 0.045824f
C17020 VDD.t1446 VSS 0.047007f
C17021 VDD.t615 VSS 0.022074f
C17022 VDD.t3260 VSS 0.020103f
C17023 VDD.t3220 VSS 0.016556f
C17024 VDD.t3259 VSS 0.035378f
C17025 VDD.t3933 VSS 0.044247f
C17026 VDD.t3931 VSS 0.021779f
C17027 VDD.t3324 VSS 0.017246f
C17028 VDD.t3322 VSS 0.023355f
C17029 VDD.t1605 VSS 0.032028f
C17030 VDD.t3504 VSS 0.025721f
C17031 VDD.t3083 VSS 0.020103f
C17032 VDD.t2222 VSS 0.034196f
C17033 VDD.t1362 VSS 0.016753f
C17034 VDD.t2 VSS 0.020103f
C17035 VDD.t3028 VSS 0.044149f
C17036 VDD.t4 VSS 0.06642f
C17037 VDD.n517 VSS 0.062606f
C17038 VDD.t362 VSS 0.02917f
C17039 VDD.t3696 VSS 0.020103f
C17040 VDD.t1468 VSS 0.021089f
C17041 VDD.t3694 VSS 0.034294f
C17042 VDD.t1765 VSS 0.024045f
C17043 VDD.t1360 VSS 0.020103f
C17044 VDD.t1430 VSS 0.025228f
C17045 VDD.t1776 VSS 0.020103f
C17046 VDD.t1467 VSS 0.020103f
C17047 VDD.t318 VSS 0.020103f
C17048 VDD.t864 VSS 0.014585f
C17049 VDD.t691 VSS 0.020498f
C17050 VDD.t17 VSS 0.030746f
C17051 VDD.t756 VSS 0.037836f
C17052 VDD.t798 VSS 0.035515f
C17053 VDD.t3505 VSS 0.019475f
C17054 VDD.t22 VSS 0.027876f
C17055 VDD.t1470 VSS 0.019475f
C17056 VDD.t1072 VSS 0.028713f
C17057 VDD.t1429 VSS 0.041166f
C17058 VDD.t3140 VSS 0.020103f
C17059 VDD.t3347 VSS 0.027002f
C17060 VDD.t741 VSS 0.031732f
C17061 VDD.t2936 VSS 0.020103f
C17062 VDD.t1352 VSS 0.02641f
C17063 VDD.t3138 VSS 0.032428f
C17064 VDD.t765 VSS 0.029816f
C17065 VDD.t3349 VSS 0.021297f
C17066 VDD.n525 VSS 0.036008f
C17067 VDD.t1894 VSS 0.023445f
C17068 VDD.t860 VSS 0.02957f
C17069 VDD.t1906 VSS 0.033015f
C17070 VDD.t61 VSS 0.037799f
C17071 VDD.t733 VSS 0.03432f
C17072 VDD.t1896 VSS 0.031982f
C17073 VDD.t3661 VSS 0.031141f
C17074 VDD.t2908 VSS 0.022074f
C17075 VDD.t3657 VSS 0.017738f
C17076 VDD.t861 VSS 0.022074f
C17077 VDD.t3659 VSS 0.024932f
C17078 VDD.t1895 VSS 0.022074f
C17079 VDD.t3663 VSS 0.020103f
C17080 VDD.t1563 VSS 0.022074f
C17081 VDD.t1592 VSS 0.028381f
C17082 VDD.t1599 VSS 0.031929f
C17083 VDD.t862 VSS 0.022074f
C17084 VDD.t1586 VSS 0.020103f
C17085 VDD.t392 VSS 0.022074f
C17086 VDD.t1597 VSS 0.036265f
C17087 VDD.t1588 VSS 0.024045f
C17088 VDD.t5 VSS 0.022074f
C17089 VDD.t779 VSS 0.042178f
C17090 VDD.t1590 VSS 0.024045f
C17091 VDD.t437 VSS 0.022074f
C17092 VDD.t1594 VSS 0.058983f
C17093 VDD.n534 VSS 0.114477f
C17094 VDD.n536 VSS 0.010255f
C17095 VDD.n542 VSS 0.010418f
C17096 VDD.n543 VSS 0.011117f
C17097 VDD.n546 VSS 0.344985f
C17098 VDD.n560 VSS 0.044473f
C17099 VDD.t396 VSS 0.050259f
C17100 VDD.t1366 VSS 0.025524f
C17101 VDD.t1705 VSS 0.027494f
C17102 VDD.t890 VSS 0.028874f
C17103 VDD.t3965 VSS 0.016556f
C17104 VDD.t892 VSS 0.020103f
C17105 VDD.t1428 VSS 0.030451f
C17106 VDD.t1364 VSS 0.03459f
C17107 VDD.t2073 VSS 0.020103f
C17108 VDD.t2505 VSS 0.016556f
C17109 VDD.t2074 VSS 0.031141f
C17110 VDD.t721 VSS 0.03252f
C17111 VDD.t3667 VSS 0.034321f
C17112 VDD.t2910 VSS 0.049197f
C17113 VDD.t1365 VSS 0.045967f
C17114 VDD.t726 VSS 0.029131f
C17115 VDD.t1427 VSS 0.031042f
C17116 VDD.t3433 VSS 0.03321f
C17117 VDD.t735 VSS 0.02444f
C17118 VDD.t744 VSS 0.024242f
C17119 VDD.t1700 VSS 0.020103f
C17120 VDD.t3375 VSS 0.038039f
C17121 VDD.n566 VSS 0.037575f
C17122 VDD.t3431 VSS 0.028184f
C17123 VDD.t2717 VSS 0.037743f
C17124 VDD.t356 VSS 0.022074f
C17125 VDD.t2713 VSS 0.020103f
C17126 VDD.t2514 VSS 0.022074f
C17127 VDD.t2715 VSS 0.033112f
C17128 VDD.t2711 VSS 0.023257f
C17129 VDD.t1611 VSS 0.021286f
C17130 VDD.t1112 VSS 0.020892f
C17131 VDD.t3901 VSS 0.020103f
C17132 VDD.t2512 VSS 0.022074f
C17133 VDD.t3895 VSS 0.020103f
C17134 VDD.t902 VSS 0.022074f
C17135 VDD.t3903 VSS 0.026805f
C17136 VDD.t3897 VSS 0.02641f
C17137 VDD.t708 VSS 0.022074f
C17138 VDD.t3909 VSS 0.034226f
C17139 VDD.t3560 VSS 0.021342f
C17140 VDD.t3905 VSS 0.026731f
C17141 VDD.t3899 VSS 0.02253f
C17142 VDD.t2513 VSS 0.02046f
C17143 VDD.t3907 VSS 0.030075f
C17144 VDD.t1111 VSS 0.028874f
C17145 VDD.t3604 VSS 0.037349f
C17146 VDD.t4024 VSS 0.02444f
C17147 VDD.t767 VSS 0.02444f
C17148 VDD.t3402 VSS 0.020103f
C17149 VDD.t1253 VSS 0.033703f
C17150 VDD.n576 VSS 0.037575f
C17151 VDD.t3602 VSS 0.028184f
C17152 VDD.t1124 VSS 0.029663f
C17153 VDD.n577 VSS 0.025355f
C17154 VDD.t1128 VSS 0.029663f
C17155 VDD.t3648 VSS 0.022074f
C17156 VDD.t1122 VSS 0.031633f
C17157 VDD.t1126 VSS 0.024735f
C17158 VDD.t1000 VSS 0.022074f
C17159 VDD.t422 VSS 0.020103f
C17160 VDD.t769 VSS 0.022074f
C17161 VDD.t432 VSS 0.02444f
C17162 VDD.t3646 VSS 0.022074f
C17163 VDD.t424 VSS 0.020103f
C17164 VDD.t3958 VSS 0.022091f
C17165 VDD.t434 VSS 0.028753f
C17166 VDD.t1568 VSS 0.021385f
C17167 VDD.t430 VSS 0.027876f
C17168 VDD.t3921 VSS 0.021385f
C17169 VDD.t426 VSS 0.029598f
C17170 VDD.t420 VSS 0.026352f
C17171 VDD.t754 VSS 0.022074f
C17172 VDD.t428 VSS 0.031141f
C17173 VDD.t1407 VSS 0.034688f
C17174 VDD.t1565 VSS 0.031535f
C17175 VDD.t1601 VSS 0.020103f
C17176 VDD.t3957 VSS 0.023651f
C17177 VDD.t3437 VSS 0.020103f
C17178 VDD.t2430 VSS 0.034491f
C17179 VDD.n586 VSS 0.037575f
C17180 VDD.t1566 VSS 0.025031f
C17181 VDD.t4123 VSS 0.023257f
C17182 VDD.t1652 VSS 0.025228f
C17183 VDD.t1658 VSS 0.044149f
C17184 VDD.t1654 VSS 0.035083f
C17185 VDD.t2974 VSS 0.022074f
C17186 VDD.t1656 VSS 0.023651f
C17187 VDD.t2768 VSS 0.022074f
C17188 VDD.t1686 VSS 0.029564f
C17189 VDD.t1694 VSS 0.033112f
C17190 VDD.t4185 VSS 0.022074f
C17191 VDD.t1690 VSS 0.022074f
C17192 VDD.t4191 VSS 0.022074f
C17193 VDD.t1696 VSS 0.022074f
C17194 VDD.t4187 VSS 0.022074f
C17195 VDD.t2601 VSS 0.022074f
C17196 VDD.t4189 VSS 0.022074f
C17197 VDD.t1688 VSS 0.022074f
C17198 VDD.t189 VSS 0.022074f
C17199 VDD.t1698 VSS 0.022074f
C17200 VDD.t201 VSS 0.022074f
C17201 VDD.t1692 VSS 0.022074f
C17202 VDD.t197 VSS 0.033112f
C17203 VDD.t193 VSS 0.035083f
C17204 VDD.t1943 VSS 0.022074f
C17205 VDD.t191 VSS 0.023651f
C17206 VDD.t1486 VSS 0.022074f
C17207 VDD.t203 VSS 0.029564f
C17208 VDD.t199 VSS 0.027002f
C17209 VDD.n600 VSS 0.025355f
C17210 VDD.t195 VSS 0.028874f
C17211 VDD.t693 VSS 0.03183f
C17212 VDD.t13 VSS 0.026312f
C17213 VDD.n601 VSS 0.037673f
C17214 VDD.t3057 VSS 0.030155f
C17215 VDD.t4125 VSS 0.022074f
C17216 VDD.t1781 VSS 0.042178f
C17217 VDD.t3059 VSS 0.034294f
C17218 VDD.t3879 VSS 0.022074f
C17219 VDD.t3061 VSS 0.020103f
C17220 VDD.t2746 VSS 0.022074f
C17221 VDD.t1384 VSS 0.020103f
C17222 VDD.t1783 VSS 0.022074f
C17223 VDD.t1378 VSS 0.020103f
C17224 VDD.t4018 VSS 0.022074f
C17225 VDD.t1372 VSS 0.031141f
C17226 VDD.t763 VSS 0.022074f
C17227 VDD.t1380 VSS 0.027313f
C17228 VDD.t1386 VSS 0.028599f
C17229 VDD.t1720 VSS 0.021385f
C17230 VDD.t1374 VSS 0.027876f
C17231 VDD.t1784 VSS 0.021385f
C17232 VDD.t1382 VSS 0.028774f
C17233 VDD.t2747 VSS 0.022106f
C17234 VDD.t1376 VSS 0.020103f
C17235 VDD.t3413 VSS 0.042276f
C17236 VDD.t736 VSS 0.031239f
C17237 VDD.n610 VSS 0.023385f
C17238 VDD.t1573 VSS 0.028184f
C17239 VDD.t2497 VSS 0.034294f
C17240 VDD.t3415 VSS 0.022074f
C17241 VDD.t2499 VSS 0.024735f
C17242 VDD.t2501 VSS 0.038039f
C17243 VDD.t2581 VSS 0.022074f
C17244 VDD.t2495 VSS 0.028184f
C17245 VDD.t239 VSS 0.033112f
C17246 VDD.t868 VSS 0.022074f
C17247 VDD.t247 VSS 0.022074f
C17248 VDD.t872 VSS 0.022074f
C17249 VDD.t243 VSS 0.022074f
C17250 VDD.t866 VSS 0.022074f
C17251 VDD.t241 VSS 0.022074f
C17252 VDD.t870 VSS 0.022074f
C17253 VDD.t249 VSS 0.022074f
C17254 VDD.t47 VSS 0.022074f
C17255 VDD.t245 VSS 0.022074f
C17256 VDD.t59 VSS 0.022074f
C17257 VDD.t273 VSS 0.022074f
C17258 VDD.t51 VSS 0.022074f
C17259 VDD.t251 VSS 0.022074f
C17260 VDD.t49 VSS 0.033112f
C17261 VDD.t55 VSS 0.038039f
C17262 VDD.t1824 VSS 0.022074f
C17263 VDD.t53 VSS 0.028184f
C17264 VDD.t45 VSS 0.044149f
C17265 VDD.t57 VSS 0.029927f
C17266 VDD.n621 VSS 0.159783f
C17267 VDD.n635 VSS 0.347695f
C17268 VDD.n636 VSS 0.302928f
C17269 VDD.n650 VSS 0.164708f
C17270 VDD.t3807 VSS 0.034667f
C17271 VDD.t3706 VSS 0.044149f
C17272 VDD.t1559 VSS 0.044149f
C17273 VDD.t1457 VSS 0.044149f
C17274 VDD.t1515 VSS 0.044149f
C17275 VDD.t1561 VSS 0.044149f
C17276 VDD.t3396 VSS 0.044149f
C17277 VDD.t3856 VSS 0.044149f
C17278 VDD.t2597 VSS 0.044149f
C17279 VDD.t2387 VSS 0.044149f
C17280 VDD.t3889 VSS 0.044149f
C17281 VDD.t3491 VSS 0.044149f
C17282 VDD.t1147 VSS 0.044149f
C17283 VDD.t4048 VSS 0.033112f
C17284 VDD.n651 VSS 0.04743f
C17285 VDD.t1293 VSS 0.066223f
C17286 VDD.n652 VSS 0.04743f
C17287 VDD.t900 VSS 0.033112f
C17288 VDD.t3210 VSS 0.044149f
C17289 VDD.t1188 VSS 0.044149f
C17290 VDD.t951 VSS 0.044149f
C17291 VDD.t3813 VSS 0.044149f
C17292 VDD.t1618 VSS 0.044149f
C17293 VDD.t2305 VSS 0.044149f
C17294 VDD.t2317 VSS 0.044149f
C17295 VDD.t3927 VSS 0.044149f
C17296 VDD.t3978 VSS 0.044149f
C17297 VDD.t4160 VSS 0.044149f
C17298 VDD.t3725 VSS 0.044149f
C17299 VDD.t949 VSS 0.044149f
C17300 VDD.t3565 VSS 0.044149f
C17301 VDD.t2155 VSS 0.044149f
C17302 VDD.t2644 VSS 0.044149f
C17303 VDD.t4015 VSS 0.033112f
C17304 VDD.t2778 VSS 0.07726f
C17305 VDD.t961 VSS 0.088298f
C17306 VDD.t3011 VSS 0.088298f
C17307 VDD.t2192 VSS 0.088298f
C17308 VDD.t986 VSS 0.088298f
C17309 VDD.t2044 VSS 0.088298f
C17310 VDD.t3563 VSS 0.07726f
C17311 VDD.n653 VSS 0.04743f
C17312 VDD.n654 VSS 0.019165f
C17313 VDD.n655 VSS 0.019165f
C17314 VDD.n656 VSS 0.019165f
C17315 VDD.n657 VSS 0.015552f
C17316 VDD.n658 VSS 0.01408f
C17317 VDD.n659 VSS 0.01013f
C17318 VDD.n675 VSS 0.011014f
C17319 VDD.n676 VSS 0.01013f
C17320 VDD.n677 VSS 0.015552f
C17321 VDD.n678 VSS 0.012957f
C17322 VDD.n680 VSS 0.378819f
C17323 VDD.n694 VSS 0.105688f
C17324 VDD.t2864 VSS 0.045006f
C17325 VDD.t1471 VSS 0.044149f
C17326 VDD.t1345 VSS 0.044149f
C17327 VDD.t4270 VSS 0.044149f
C17328 VDD.t1900 VSS 0.044149f
C17329 VDD.t2831 VSS 0.044149f
C17330 VDD.t4005 VSS 0.044149f
C17331 VDD.t1557 VSS 0.044149f
C17332 VDD.t3673 VSS 0.044149f
C17333 VDD.t3119 VSS 0.044149f
C17334 VDD.t2821 VSS 0.044149f
C17335 VDD.t3371 VSS 0.044149f
C17336 VDD.t1321 VSS 0.044149f
C17337 VDD.t1186 VSS 0.044149f
C17338 VDD.t3708 VSS 0.069504f
C17339 VDD.t3867 VSS 0.044149f
C17340 VDD.t2849 VSS 0.044149f
C17341 VDD.t2958 VSS 0.044149f
C17342 VDD.t2414 VSS 0.044149f
C17343 VDD.t918 VSS 0.044149f
C17344 VDD.t3712 VSS 0.044149f
C17345 VDD.t927 VSS 0.044149f
C17346 VDD.t935 VSS 0.044149f
C17347 VDD.t2979 VSS 0.044149f
C17348 VDD.t1498 VSS 0.044149f
C17349 VDD.t1343 VSS 0.044149f
C17350 VDD.t3441 VSS 0.044149f
C17351 VDD.t2579 VSS 0.044149f
C17352 VDD.t3593 VSS 0.044149f
C17353 VDD.t3917 VSS 0.044149f
C17354 VDD.t1136 VSS 0.044149f
C17355 VDD.t3935 VSS 0.044149f
C17356 VDD.t1793 VSS 0.044149f
C17357 VDD.t2491 VSS 0.044149f
C17358 VDD.t1437 VSS 0.044149f
C17359 VDD.t3367 VSS 0.044149f
C17360 VDD.t3164 VSS 0.044149f
C17361 VDD.t1149 VSS 0.044149f
C17362 VDD.t2845 VSS 0.044149f
C17363 VDD.t4143 VSS 0.044149f
C17364 VDD.t3160 VSS 0.044149f
C17365 VDD.t2966 VSS 0.044149f
C17366 VDD.t2216 VSS 0.044149f
C17367 VDD.t2833 VSS 0.044149f
C17368 VDD.t1539 VSS 0.044149f
C17369 VDD.t2404 VSS 0.044149f
C17370 VDD.t1979 VSS 0.044149f
C17371 VDD.t3439 VSS 0.069504f
C17372 VDD.n706 VSS 0.012547f
C17373 VDD.n707 VSS 0.01013f
C17374 VDD.n724 VSS 0.012547f
C17375 VDD.n727 VSS 0.118404f
C17376 VDD.n741 VSS 0.105688f
C17377 VDD.t3449 VSS 0.045006f
C17378 VDD.t3423 VSS 0.044149f
C17379 VDD.t3805 VSS 0.044149f
C17380 VDD.t1332 VSS 0.044149f
C17381 VDD.t3642 VSS 0.044149f
C17382 VDD.t3963 VSS 0.044149f
C17383 VDD.t4163 VSS 0.044149f
C17384 VDD.t1616 VSS 0.044149f
C17385 VDD.t4156 VSS 0.044149f
C17386 VDD.t3995 VSS 0.044149f
C17387 VDD.t1224 VSS 0.044149f
C17388 VDD.t3041 VSS 0.044149f
C17389 VDD.t3110 VSS 0.044149f
C17390 VDD.t4225 VSS 0.044149f
C17391 VDD.t2255 VSS 0.069504f
C17392 VDD.t2275 VSS 0.044149f
C17393 VDD.t4150 VSS 0.044149f
C17394 VDD.t1761 VSS 0.044149f
C17395 VDD.t1097 VSS 0.044149f
C17396 VDD.t1289 VSS 0.044149f
C17397 VDD.t1417 VSS 0.044149f
C17398 VDD.t2944 VSS 0.044149f
C17399 VDD.t1832 VSS 0.044149f
C17400 VDD.t2297 VSS 0.044149f
C17401 VDD.t2372 VSS 0.044149f
C17402 VDD.t3178 VSS 0.044149f
C17403 VDD.t933 VSS 0.044149f
C17404 VDD.t3636 VSS 0.044149f
C17405 VDD.t1247 VSS 0.044149f
C17406 VDD.t1179 VSS 0.044149f
C17407 VDD.t2063 VSS 0.044149f
C17408 VDD.t4272 VSS 0.069504f
C17409 VDD.t1249 VSS 0.044149f
C17410 VDD.t2652 VSS 0.044149f
C17411 VDD.t2207 VSS 0.044149f
C17412 VDD.t1421 VSS 0.044149f
C17413 VDD.t1388 VSS 0.044149f
C17414 VDD.t2485 VSS 0.044149f
C17415 VDD.t1674 VSS 0.044149f
C17416 VDD.t2991 VSS 0.044149f
C17417 VDD.t3373 VSS 0.044149f
C17418 VDD.t3971 VSS 0.044149f
C17419 VDD.t2703 VSS 0.044149f
C17420 VDD.t1724 VSS 0.044149f
C17421 VDD.t2603 VSS 0.044149f
C17422 VDD.t3427 VSS 0.044149f
C17423 VDD.t2422 VSS 0.044149f
C17424 VDD.t2872 VSS 0.044149f
C17425 VDD.t1785 VSS 0.069504f
C17426 VDD.t4103 VSS 0.044149f
C17427 VDD.t2533 VSS 0.044149f
C17428 VDD.t3158 VSS 0.044149f
C17429 VDD.t1975 VSS 0.044149f
C17430 VDD.t3671 VSS 0.044149f
C17431 VDD.t3455 VSS 0.044149f
C17432 VDD.t2575 VSS 0.044149f
C17433 VDD.t1433 VSS 0.044149f
C17434 VDD.t3435 VSS 0.044149f
C17435 VDD.t3404 VSS 0.044149f
C17436 VDD.t3266 VSS 0.044149f
C17437 VDD.t2537 VSS 0.044149f
C17438 VDD.t3584 VSS 0.044149f
C17439 VDD.t3484 VSS 0.044149f
C17440 VDD.t3034 VSS 0.044149f
C17441 VDD.t3787 VSS 0.044149f
C17442 VDD.t1337 VSS 0.040207f
C17443 VDD.t643 VSS 0.044149f
C17444 VDD.t3520 VSS 0.052033f
C17445 VDD.t19 VSS 0.044149f
C17446 VDD.t3679 VSS 0.02917f
C17447 VDD.t959 VSS 0.044149f
C17448 VDD.t3379 VSS 0.044149f
C17449 VDD.t4203 VSS 0.044149f
C17450 VDD.t3937 VSS 0.044149f
C17451 VDD.t3100 VSS 0.044149f
C17452 VDD.t923 VSS 0.044149f
C17453 VDD.t2815 VSS 0.044149f
C17454 VDD.t3809 VSS 0.044149f
C17455 VDD.t3240 VSS 0.044149f
C17456 VDD.t1241 VSS 0.044149f
C17457 VDD.t914 VSS 0.055186f
C17458 VDD.t931 VSS 0.080541f
C17459 VDD.n748 VSS 0.01408f
C17460 VDD.n749 VSS 0.01013f
C17461 VDD.n766 VSS 0.012547f
C17462 VDD.n767 VSS 0.01013f
C17463 VDD.n785 VSS 0.012547f
C17464 VDD.n786 VSS 0.01013f
C17465 VDD.n803 VSS 0.012547f
C17466 VDD.n806 VSS 0.118404f
C17467 VDD.n820 VSS 0.105688f
C17468 VDD.t2007 VSS 0.045006f
C17469 VDD.t2829 VSS 0.044149f
C17470 VDD.t2209 VSS 0.044149f
C17471 VDD.t2661 VSS 0.044149f
C17472 VDD.t2159 VSS 0.044149f
C17473 VDD.t4286 VSS 0.044149f
C17474 VDD.t4280 VSS 0.044149f
C17475 VDD.t2902 VSS 0.044149f
C17476 VDD.t1099 VSS 0.044149f
C17477 VDD.t3102 VSS 0.044149f
C17478 VDD.t4076 VSS 0.044149f
C17479 VDD.t2398 VSS 0.044149f
C17480 VDD.t2448 VSS 0.044149f
C17481 VDD.t2303 VSS 0.044149f
C17482 VDD.t3156 VSS 0.069504f
C17483 VDD.t3236 VSS 0.044149f
C17484 VDD.t3881 VSS 0.044149f
C17485 VDD.t1632 VSS 0.044149f
C17486 VDD.t2839 VSS 0.044149f
C17487 VDD.t1684 VSS 0.044149f
C17488 VDD.t4101 VSS 0.044149f
C17489 VDD.t3842 VSS 0.044149f
C17490 VDD.t1982 VSS 0.044149f
C17491 VDD.t3003 VSS 0.044149f
C17492 VDD.t2954 VSS 0.044149f
C17493 VDD.t3277 VSS 0.044149f
C17494 VDD.t1350 VSS 0.044149f
C17495 VDD.t1802 VSS 0.044149f
C17496 VDD.t3005 VSS 0.044149f
C17497 VDD.t2900 VSS 0.044149f
C17498 VDD.t3425 VSS 0.044149f
C17499 VDD.t1190 VSS 0.044149f
C17500 VDD.t4158 VSS 0.044149f
C17501 VDD.t3013 VSS 0.044149f
C17502 VDD.t4292 VSS 0.044149f
C17503 VDD.t2462 VSS 0.044149f
C17504 VDD.t3477 VSS 0.044149f
C17505 VDD.t2402 VSS 0.044149f
C17506 VDD.t971 VSS 0.044149f
C17507 VDD.t3718 VSS 0.044149f
C17508 VDD.t4169 VSS 0.044149f
C17509 VDD.t3654 VSS 0.044149f
C17510 VDD.t2042 VSS 0.044149f
C17511 VDD.t4218 VSS 0.044149f
C17512 VDD.t1990 VSS 0.044149f
C17513 VDD.t2476 VSS 0.044149f
C17514 VDD.t3152 VSS 0.044149f
C17515 VDD.t3783 VSS 0.069504f
C17516 VDD.n832 VSS 0.012547f
C17517 VDD.n833 VSS 0.01013f
C17518 VDD.n850 VSS 0.012547f
C17519 VDD.n853 VSS 0.118404f
C17520 VDD.n867 VSS 0.105688f
C17521 VDD.t3049 VSS 0.045006f
C17522 VDD.t1739 VSS 0.044149f
C17523 VDD.t3469 VSS 0.044149f
C17524 VDD.t3640 VSS 0.044149f
C17525 VDD.t2157 VSS 0.044149f
C17526 VDD.t3923 VSS 0.044149f
C17527 VDD.t4177 VSS 0.044149f
C17528 VDD.t1259 VSS 0.044149f
C17529 VDD.t4171 VSS 0.044149f
C17530 VDD.t2560 VSS 0.044149f
C17531 VDD.t1226 VSS 0.044149f
C17532 VDD.t3665 VSS 0.044149f
C17533 VDD.t3112 VSS 0.044149f
C17534 VDD.t4227 VSS 0.044149f
C17535 VDD.t2315 VSS 0.069504f
C17536 VDD.t2125 VSS 0.044149f
C17537 VDD.t4167 VSS 0.044149f
C17538 VDD.t3381 VSS 0.044149f
C17539 VDD.t1245 VSS 0.044149f
C17540 VDD.t3688 VSS 0.044149f
C17541 VDD.t1228 VSS 0.044149f
C17542 VDD.t3536 VSS 0.044149f
C17543 VDD.t4011 VSS 0.044149f
C17544 VDD.t2721 VSS 0.044149f
C17545 VDD.t2642 VSS 0.044149f
C17546 VDD.t3451 VSS 0.044149f
C17547 VDD.t1297 VSS 0.044149f
C17548 VDD.t3345 VSS 0.044149f
C17549 VDD.t1251 VSS 0.044149f
C17550 VDD.t3091 VSS 0.044149f
C17551 VDD.t2172 VSS 0.044149f
C17552 VDD.t3136 VSS 0.044149f
C17553 VDD.t2520 VSS 0.044149f
C17554 VDD.t1737 VSS 0.044149f
C17555 VDD.t2640 VSS 0.044149f
C17556 VDD.t1732 VSS 0.044149f
C17557 VDD.t3252 VSS 0.044149f
C17558 VDD.t3999 VSS 0.044149f
C17559 VDD.t3377 VSS 0.044149f
C17560 VDD.t3929 VSS 0.044149f
C17561 VDD.t3528 VSS 0.044149f
C17562 VDD.t965 VSS 0.044149f
C17563 VDD.t939 VSS 0.044149f
C17564 VDD.t3976 VSS 0.044149f
C17565 VDD.t1195 VSS 0.044149f
C17566 VDD.t1679 VSS 0.044149f
C17567 VDD.t1370 VSS 0.044149f
C17568 VDD.t2526 VSS 0.069504f
C17569 VDD.n879 VSS 0.012547f
C17570 VDD.n880 VSS 0.01013f
C17571 VDD.n897 VSS 0.012547f
C17572 VDD.n900 VSS 0.118404f
C17573 VDD.n914 VSS 0.105688f
C17574 VDD.t3419 VSS 0.045006f
C17575 VDD.t3591 VSS 0.044149f
C17576 VDD.t4207 VSS 0.044149f
C17577 VDD.t1134 VSS 0.044149f
C17578 VDD.t1481 VSS 0.044149f
C17579 VDD.t3074 VSS 0.044149f
C17580 VDD.t2800 VSS 0.044149f
C17581 VDD.t1582 VSS 0.044149f
C17582 VDD.t4201 VSS 0.044149f
C17583 VDD.t1138 VSS 0.044149f
C17584 VDD.t898 VSS 0.044149f
C17585 VDD.t2725 VSS 0.044149f
C17586 VDD.t4213 VSS 0.044149f
C17587 VDD.t3081 VSS 0.044149f
C17588 VDD.t2940 VSS 0.069504f
C17589 VDD.t3941 VSS 0.044149f
C17590 VDD.t1620 VSS 0.044149f
C17591 VDD.t3318 VSS 0.044149f
C17592 VDD.t3947 VSS 0.044149f
C17593 VDD.t2843 VSS 0.044149f
C17594 VDD.t2420 VSS 0.044149f
C17595 VDD.t1212 VSS 0.044149f
C17596 VDD.t1423 VSS 0.044149f
C17597 VDD.t3988 VSS 0.044149f
C17598 VDD.t1535 VSS 0.044149f
C17599 VDD.t1707 VSS 0.044149f
C17600 VDD.t1937 VSS 0.044149f
C17601 VDD.t3838 VSS 0.044149f
C17602 VDD.t3162 VSS 0.044149f
C17603 VDD.t3238 VSS 0.044149f
C17604 VDD.t2092 VSS 0.044149f
C17605 VDD.t3043 VSS 0.080541f
C17606 VDD.t2707 VSS 0.055186f
C17607 VDD.t2201 VSS 0.044149f
C17608 VDD.t4238 VSS 0.044149f
C17609 VDD.t3832 VSS 0.044149f
C17610 VDD.t2823 VSS 0.044149f
C17611 VDD.t1889 VSS 0.044149f
C17612 VDD.t2301 VSS 0.044149f
C17613 VDD.t3421 VSS 0.044149f
C17614 VDD.t3187 VSS 0.044149f
C17615 VDD.t2084 VSS 0.044149f
C17616 VDD.t3290 VSS 0.044149f
C17617 VDD.t4232 VSS 0.044149f
C17618 VDD.t1730 VSS 0.044149f
C17619 VDD.t984 VSS 0.044149f
C17620 VDD.t2835 VSS 0.044149f
C17621 VDD.t3684 VSS 0.033112f
C17622 VDD.n915 VSS 0.04743f
C17623 VDD.t3457 VSS 0.033112f
C17624 VDD.t2029 VSS 0.044149f
C17625 VDD.t2061 VSS 0.044149f
C17626 VDD.t3369 VSS 0.044149f
C17627 VDD.t1777 VSS 0.044149f
C17628 VDD.t1984 VSS 0.044149f
C17629 VDD.t1479 VSS 0.044149f
C17630 VDD.t2554 VSS 0.044149f
C17631 VDD.t3015 VSS 0.037053f
C17632 VDD.t4064 VSS 0.044149f
C17633 VDD.t2295 VSS 0.048288f
C17634 VDD.t3534 VSS 0.040601f
C17635 VDD.t3077 VSS 0.036068f
C17636 VDD.t2432 VSS 0.016556f
C17637 VDD.t3076 VSS 0.041192f
C17638 VDD.t2313 VSS 0.042966f
C17639 VDD.t2859 VSS 0.02444f
C17640 VDD.t3329 VSS 0.016556f
C17641 VDD.t2857 VSS 0.033703f
C17642 VDD.t2083 VSS 0.025819f
C17643 VDD.t1672 VSS 0.025228f
C17644 VDD.t3753 VSS 0.030746f
C17645 VDD.t236 VSS 0.02917f
C17646 VDD.t1506 VSS 0.023651f
C17647 VDD.t2620 VSS 0.022074f
C17648 VDD.t645 VSS 0.024045f
C17649 VDD.t3982 VSS 0.039221f
C17650 VDD.t4300 VSS 0.037743f
C17651 VDD.t1512 VSS 0.02917f
C17652 VDD.t636 VSS 0.020103f
C17653 VDD.t897 VSS 0.031633f
C17654 VDD.t3722 VSS 0.040207f
C17655 VDD.t2412 VSS 0.037842f
C17656 VDD.t3355 VSS 0.035575f
C17657 VDD.t1834 VSS 0.03252f
C17658 VDD.t4297 VSS 0.031239f
C17659 VDD.t4299 VSS 0.034393f
C17660 VDD.t2088 VSS 0.039911f
C17661 VDD.t3703 VSS 0.0271f
C17662 VDD.t877 VSS 0.016556f
C17663 VDD.t3705 VSS 0.016556f
C17664 VDD.t878 VSS 0.0271f
C17665 VDD.t2309 VSS 0.03794f
C17666 VDD.t3186 VSS 0.032422f
C17667 VDD.t3184 VSS 0.017738f
C17668 VDD.n919 VSS 0.031268f
C17669 VDD.n923 VSS 0.010974f
C17670 VDD.n924 VSS 0.014938f
C17671 VDD.n925 VSS 0.013432f
C17672 VDD.n926 VSS 0.015243f
C17673 VDD.n928 VSS 0.015958f
C17674 VDD.n929 VSS 0.011166f
C17675 VDD.n931 VSS 0.015714f
C17676 VDD.n932 VSS 0.014181f
C17677 VDD.n941 VSS 0.01408f
C17678 VDD.n942 VSS 0.01013f
C17679 VDD.n959 VSS 0.01408f
C17680 VDD.n960 VSS 0.01013f
C17681 VDD.n977 VSS 0.012547f
C17682 VDD.n980 VSS 0.118404f
C17683 VDD.n994 VSS 0.105688f
C17684 VDD.t2798 VSS 0.045006f
C17685 VDD.t3745 VSS 0.044149f
C17686 VDD.t1789 VSS 0.044149f
C17687 VDD.t2962 VSS 0.044149f
C17688 VDD.t2729 VSS 0.044149f
C17689 VDD.t2870 VSS 0.044149f
C17690 VDD.t2896 VSS 0.044149f
C17691 VDD.t1510 VSS 0.044149f
C17692 VDD.t2214 VSS 0.044149f
C17693 VDD.t2038 VSS 0.044149f
C17694 VDD.t2667 VSS 0.044149f
C17695 VDD.t3893 VSS 0.044149f
C17696 VDD.t977 VSS 0.044149f
C17697 VDD.t1628 VSS 0.044149f
C17698 VDD.t2774 VSS 0.069504f
C17699 VDD.t4038 VSS 0.044149f
C17700 VDD.t3198 VSS 0.044149f
C17701 VDD.t2368 VSS 0.044149f
C17702 VDD.t2361 VSS 0.044149f
C17703 VDD.t2251 VSS 0.044149f
C17704 VDD.t2669 VSS 0.044149f
C17705 VDD.t2253 VSS 0.044149f
C17706 VDD.t3949 VSS 0.044149f
C17707 VDD.t1682 VSS 0.044149f
C17708 VDD.t4042 VSS 0.044149f
C17709 VDD.t2860 VSS 0.044149f
C17710 VDD.t4096 VSS 0.044149f
C17711 VDD.t1231 VSS 0.044149f
C17712 VDD.t2489 VSS 0.044149f
C17713 VDD.t3279 VSS 0.044149f
C17714 VDD.t3686 VSS 0.044149f
C17715 VDD.t1810 VSS 0.044149f
C17716 VDD.t3586 VSS 0.044149f
C17717 VDD.t2807 VSS 0.044149f
C17718 VDD.t1718 VSS 0.044149f
C17719 VDD.t3986 VSS 0.044149f
C17720 VDD.t2450 VSS 0.044149f
C17721 VDD.t3087 VSS 0.044149f
C17722 VDD.t2277 VSS 0.044149f
C17723 VDD.t2101 VSS 0.044149f
C17724 VDD.t4199 VSS 0.044149f
C17725 VDD.t1812 VSS 0.044149f
C17726 VDD.t3572 VSS 0.044149f
C17727 VDD.t3574 VSS 0.044149f
C17728 VDD.t2757 VSS 0.044149f
C17729 VDD.t1800 VSS 0.044149f
C17730 VDD.t2493 VSS 0.044149f
C17731 VDD.t1439 VSS 0.069504f
C17732 VDD.n1006 VSS 0.012547f
C17733 VDD.n1007 VSS 0.01013f
C17734 VDD.n1024 VSS 0.012547f
C17735 VDD.n1027 VSS 0.118404f
C17736 VDD.n1041 VSS 0.105688f
C17737 VDD.t4282 VSS 0.045006f
C17738 VDD.t3803 VSS 0.044149f
C17739 VDD.t3799 VSS 0.044149f
C17740 VDD.t2119 VSS 0.044149f
C17741 VDD.t1914 VSS 0.044149f
C17742 VDD.t2027 VSS 0.044149f
C17743 VDD.t4276 VSS 0.044149f
C17744 VDD.t3248 VSS 0.044149f
C17745 VDD.t998 VSS 0.044149f
C17746 VDD.t2868 VSS 0.044149f
C17747 VDD.t3567 VSS 0.044149f
C17748 VDD.t1291 VSS 0.044149f
C17749 VDD.t4040 VSS 0.044149f
C17750 VDD.t3576 VSS 0.044149f
C17751 VDD.t2583 VSS 0.069504f
C17752 VDD.t2330 VSS 0.044149f
C17753 VDD.t1865 VSS 0.044149f
C17754 VDD.t3007 VSS 0.044149f
C17755 VDD.t2675 VSS 0.044149f
C17756 VDD.t3682 VSS 0.044149f
C17757 VDD.t3154 VSS 0.044149f
C17758 VDD.t3108 VSS 0.044149f
C17759 VDD.t3515 VSS 0.044149f
C17760 VDD.t975 VSS 0.044149f
C17761 VDD.t3353 VSS 0.044149f
C17762 VDD.t2359 VSS 0.044149f
C17763 VDD.t1409 VSS 0.044149f
C17764 VDD.t3142 VSS 0.044149f
C17765 VDD.t2659 VSS 0.044149f
C17766 VDD.t4068 VSS 0.044149f
C17767 VDD.t3751 VSS 0.044149f
C17768 VDD.t3311 VSS 0.044149f
C17769 VDD.t2809 VSS 0.044149f
C17770 VDD.t2590 VSS 0.044149f
C17771 VDD.t3384 VSS 0.044149f
C17772 VDD.t1233 VSS 0.044149f
C17773 VDD.t4197 VSS 0.044149f
C17774 VDD.t1910 VSS 0.044149f
C17775 VDD.t3885 VSS 0.044149f
C17776 VDD.t1415 VSS 0.044149f
C17777 VDD.t3262 VSS 0.044149f
C17778 VDD.t3853 VSS 0.044149f
C17779 VDD.t3634 VSS 0.044149f
C17780 VDD.t2299 VSS 0.044149f
C17781 VDD.t2546 VSS 0.044149f
C17782 VDD.t3522 VSS 0.044149f
C17783 VDD.t2127 VSS 0.044149f
C17784 VDD.t1130 VSS 0.069504f
C17785 VDD.n1053 VSS 0.012547f
C17786 VDD.n1054 VSS 0.01013f
C17787 VDD.n1071 VSS 0.012547f
C17788 VDD.n1074 VSS 0.118404f
C17789 VDD.n1088 VSS 0.105688f
C17790 VDD.t2522 VSS 0.045006f
C17791 VDD.t1626 VSS 0.044149f
C17792 VDD.t2291 VSS 0.044149f
C17793 VDD.t2912 VSS 0.044149f
C17794 VDD.t2380 VSS 0.044149f
C17795 VDD.t2031 VSS 0.044149f
C17796 VDD.t3341 VSS 0.044149f
C17797 VDD.t1912 VSS 0.044149f
C17798 VDD.t3117 VSS 0.044149f
C17799 VDD.t1922 VSS 0.044149f
C17800 VDD.t3453 VSS 0.044149f
C17801 VDD.t3939 VSS 0.044149f
C17802 VDD.t1411 VSS 0.044149f
C17803 VDD.t1722 VSS 0.044149f
C17804 VDD.t967 VSS 0.069504f
C17805 VDD.t2898 VSS 0.044149f
C17806 VDD.t1443 VSS 0.044149f
C17807 VDD.t4020 VSS 0.044149f
C17808 VDD.t1857 VSS 0.044149f
C17809 VDD.t1992 VSS 0.044149f
C17810 VDD.t2036 VSS 0.044149f
C17811 VDD.t1339 VSS 0.044149f
C17812 VDD.t4183 VSS 0.044149f
C17813 VDD.t2321 VSS 0.044149f
C17814 VDD.t4105 VSS 0.044149f
C17815 VDD.t2942 VSS 0.044149f
C17816 VDD.t4053 VSS 0.044149f
C17817 VDD.t3398 VSS 0.044149f
C17818 VDD.t1840 VSS 0.044149f
C17819 VDD.t3070 VSS 0.044149f
C17820 VDD.t3811 VSS 0.044149f
C17821 VDD.t4181 VSS 0.080541f
C17822 VDD.t2677 VSS 0.055186f
C17823 VDD.t2665 VSS 0.044149f
C17824 VDD.t3524 VSS 0.044149f
C17825 VDD.t2790 VSS 0.044149f
C17826 VDD.t3967 VSS 0.044149f
C17827 VDD.t2874 VSS 0.044149f
C17828 VDD.t3129 VSS 0.044149f
C17829 VDD.t4072 VSS 0.044149f
C17830 VDD.t2444 VSS 0.044149f
C17831 VDD.t1358 VSS 0.044149f
C17832 VDD.t1523 VSS 0.044149f
C17833 VDD.t2269 VSS 0.044149f
C17834 VDD.t3406 VSS 0.044149f
C17835 VDD.t1235 VSS 0.044149f
C17836 VDD.t2112 VSS 0.044149f
C17837 VDD.t4066 VSS 0.033112f
C17838 VDD.n1089 VSS 0.04743f
C17839 VDD.t1243 VSS 0.026016f
C17840 VDD.t480 VSS 0.044149f
C17841 VDD.t2393 VSS 0.044149f
C17842 VDD.t4121 VSS 0.039221f
C17843 VDD.t443 VSS 0.044149f
C17844 VDD.t758 VSS 0.024045f
C17845 VDD.t815 VSS 0.03528f
C17846 VDD.t823 VSS 0.031239f
C17847 VDD.t4115 VSS 0.024045f
C17848 VDD.t445 VSS 0.020103f
C17849 VDD.t3755 VSS 0.023651f
C17850 VDD.t289 VSS 0.036955f
C17851 VDD.t283 VSS 0.024045f
C17852 VDD.t297 VSS 0.020103f
C17853 VDD.t1284 VSS 0.020103f
C17854 VDD.t291 VSS 0.027593f
C17855 VDD.t293 VSS 0.030746f
C17856 VDD.t1255 VSS 0.020103f
C17857 VDD.t285 VSS 0.020103f
C17858 VDD.t4261 VSS 0.024045f
C17859 VDD.t295 VSS 0.020103f
C17860 VDD.t1286 VSS 0.020103f
C17861 VDD.t299 VSS 0.020103f
C17862 VDD.t2751 VSS 0.024045f
C17863 VDD.t287 VSS 0.031141f
C17864 VDD.t751 VSS 0.03252f
C17865 VDD.t2532 VSS 0.033799f
C17866 VDD.t1033 VSS 0.024045f
C17867 VDD.t3096 VSS 0.020103f
C17868 VDD.t1220 VSS 0.029958f
C17869 VDD.t1035 VSS 0.034688f
C17870 VDD.t2268 VSS 0.039419f
C17871 VDD.t916 VSS 0.025228f
C17872 VDD.t1295 VSS 0.023651f
C17873 VDD.t3630 VSS 0.024045f
C17874 VDD.t3064 VSS 0.027396f
C17875 VDD.t3066 VSS 0.038532f
C17876 VDD.t880 VSS 0.049963f
C17877 VDD.t3973 VSS 0.041389f
C17878 VDD.t4175 VSS 0.016556f
C17879 VDD.t3975 VSS 0.034294f
C17880 VDD.t1550 VSS 0.044937f
C17881 VDD.t1556 VSS 0.020103f
C17882 VDD.t727 VSS 0.016556f
C17883 VDD.t1554 VSS 0.02444f
C17884 VDD.t4173 VSS 0.022074f
C17885 VDD.t2528 VSS 0.020103f
C17886 VDD.t4260 VSS 0.018724f
C17887 VDD.t1197 VSS 0.041028f
C17888 VDD.t848 VSS 0.043887f
C17889 VDD.n1097 VSS 0.039013f
C17890 VDD.n1098 VSS 0.027523f
C17891 VDD.n1101 VSS 0.010742f
C17892 VDD.n1103 VSS 0.013035f
C17893 VDD.n1104 VSS 0.015445f
C17894 VDD.n1106 VSS 0.011288f
C17895 VDD.n1109 VSS 0.011083f
C17896 VDD.n1118 VSS 0.013761f
C17897 VDD.n1119 VSS 0.015714f
C17898 VDD.n1120 VSS 0.010568f
C17899 VDD.n1121 VSS 0.01408f
C17900 VDD.n1122 VSS 0.01013f
C17901 VDD.n1139 VSS 0.01408f
C17902 VDD.n1140 VSS 0.01013f
C17903 VDD.n1157 VSS 0.012547f
C17904 VDD.n1160 VSS 0.118404f
C17905 VDD.n1174 VSS 0.105688f
C17906 VDD.t4290 VSS 0.045006f
C17907 VDD.t3789 VSS 0.044149f
C17908 VDD.t3173 VSS 0.044149f
C17909 VDD.t4211 VSS 0.044149f
C17910 VDD.t3246 VSS 0.044149f
C17911 VDD.t1473 VSS 0.044149f
C17912 VDD.t1354 VSS 0.044149f
C17913 VDD.t4266 VSS 0.044149f
C17914 VDD.t2013 VSS 0.044149f
C17915 VDD.t1207 VSS 0.044149f
C17916 VDD.t2483 VSS 0.044149f
C17917 VDD.t3250 VSS 0.044149f
C17918 VDD.t2395 VSS 0.044149f
C17919 VDD.t3132 VSS 0.044149f
C17920 VDD.t3001 VSS 0.080541f
C17921 VDD.t3098 VSS 0.066223f
C17922 VDD.t3969 VSS 0.044149f
C17923 VDD.t3883 VSS 0.044149f
C17924 VDD.t3556 VSS 0.044149f
C17925 VDD.t2446 VSS 0.044149f
C17926 VDD.t3549 VSS 0.044149f
C17927 VDD.t3134 VSS 0.044149f
C17928 VDD.t1630 VSS 0.044149f
C17929 VDD.t2418 VSS 0.044149f
C17930 VDD.t2123 VSS 0.044149f
C17931 VDD.t1299 VSS 0.044149f
C17932 VDD.t2701 VSS 0.044149f
C17933 VDD.t2552 VSS 0.044149f
C17934 VDD.t990 VSS 0.044149f
C17935 VDD.t2106 VSS 0.044149f
C17936 VDD.t3764 VSS 0.033112f
C17937 VDD.t1816 VSS 0.027002f
C17938 VDD.t1814 VSS 0.028184f
C17939 VDD.t2573 VSS 0.022074f
C17940 VDD.t1818 VSS 0.038039f
C17941 VDD.t1996 VSS 0.028184f
C17942 VDD.t1451 VSS 0.022074f
C17943 VDD.t1820 VSS 0.038039f
C17944 VDD.t1994 VSS 0.038532f
C17945 VDD.t1199 VSS 0.022074f
C17946 VDD.t1822 VSS 0.027691f
C17947 VDD.t1999 VSS 0.026903f
C17948 VDD.t2163 VSS 0.021385f
C17949 VDD.t2165 VSS 0.041488f
C17950 VDD.t1998 VSS 0.044937f
C17951 VDD.t1146 VSS 0.036561f
C17952 VDD.t1144 VSS 0.017049f
C17953 VDD.t2647 VSS 0.022074f
C17954 VDD.t846 VSS 0.044149f
C17955 VDD.t2178 VSS 0.044641f
C17956 VDD.t3945 VSS 0.044149f
C17957 VDD.t3009 VSS 0.044149f
C17958 VDD.t969 VSS 0.055186f
C17959 VDD.n1175 VSS 0.04743f
C17960 VDD.n1179 VSS 0.015404f
C17961 VDD.n1180 VSS 0.013295f
C17962 VDD.n1181 VSS 0.010061f
C17963 VDD.n1182 VSS 0.012648f
C17964 VDD.n1186 VSS 0.01408f
C17965 VDD.n1187 VSS 0.01013f
C17966 VDD.n1202 VSS 0.010568f
C17967 VDD.n1203 VSS 0.01408f
C17968 VDD.n1206 VSS 0.118404f
C17969 VDD.n1220 VSS 0.105688f
C17970 VDD.t2249 VSS 0.045006f
C17971 VDD.t2151 VSS 0.044149f
C17972 VDD.t2182 VSS 0.044149f
C17973 VDD.t3747 VSS 0.044149f
C17974 VDD.t2391 VSS 0.044149f
C17975 VDD.t2129 VSS 0.044149f
C17976 VDD.t2134 VSS 0.044149f
C17977 VDD.t2363 VSS 0.044149f
C17978 VDD.t2888 VSS 0.044149f
C17979 VDD.t3821 VSS 0.044149f
C17980 VDD.t1986 VSS 0.044149f
C17981 VDD.t3915 VSS 0.044149f
C17982 VDD.t3202 VSS 0.044149f
C17983 VDD.t3846 VSS 0.044149f
C17984 VDD.t893 VSS 0.069504f
C17985 VDD.t3531 VSS 0.044149f
C17986 VDD.t1500 VSS 0.044149f
C17987 VDD.t3417 VSS 0.044149f
C17988 VDD.t957 VSS 0.044149f
C17989 VDD.t3873 VSS 0.044149f
C17990 VDD.t2709 VSS 0.044149f
C17991 VDD.t3913 VSS 0.044149f
C17992 VDD.t3793 VSS 0.044149f
C17993 VDD.t2673 VSS 0.044149f
C17994 VDD.t2539 VSS 0.044149f
C17995 VDD.t2071 VSS 0.044149f
C17996 VDD.t1431 VSS 0.044149f
C17997 VDD.t1537 VSS 0.044149f
C17998 VDD.t2934 VSS 0.044149f
C17999 VDD.t1116 VSS 0.044149f
C18000 VDD.t2558 VSS 0.044149f
C18001 VDD.t4082 VSS 0.033703f
C18002 VDD.t4080 VSS 0.028381f
C18003 VDD.t2326 VSS 0.020103f
C18004 VDD.t4088 VSS 0.039813f
C18005 VDD.t4084 VSS 0.028381f
C18006 VDD.t2993 VSS 0.043557f
C18007 VDD.t4033 VSS 0.046317f
C18008 VDD.t703 VSS 0.044149f
C18009 VDD.t3610 VSS 0.044149f
C18010 VDD.t324 VSS 0.044149f
C18011 VDD.t2794 VSS 0.081202f
C18012 VDD.t2228 VSS 0.088298f
C18013 VDD.t1546 VSS 0.088298f
C18014 VDD.t1455 VSS 0.088298f
C18015 VDD.t3614 VSS 0.080541f
C18016 VDD.n1221 VSS 0.015714f
C18017 VDD.n1222 VSS 0.019165f
C18018 VDD.n1223 VSS 0.019165f
C18019 VDD.n1224 VSS 0.019165f
C18020 VDD.n1225 VSS 0.017084f
C18021 VDD.n1226 VSS 0.01408f
C18022 VDD.n1227 VSS 0.01013f
C18023 VDD.n1244 VSS 0.012547f
C18024 VDD.n1247 VSS 0.118404f
C18025 VDD.n1261 VSS 0.105688f
C18026 VDD.t4294 VSS 0.045006f
C18027 VDD.t2759 VSS 0.044149f
C18028 VDD.t3206 VSS 0.044149f
C18029 VDD.t3578 VSS 0.044149f
C18030 VDD.t3045 VSS 0.044149f
C18031 VDD.t2780 VSS 0.044149f
C18032 VDD.t3836 VSS 0.044149f
C18033 VDD.t982 VSS 0.044149f
C18034 VDD.t3464 VSS 0.044149f
C18035 VDD.t1214 VSS 0.044149f
C18036 VDD.t1580 VSS 0.044149f
C18037 VDD.t2025 VSS 0.044149f
C18038 VDD.t2681 VSS 0.044149f
C18039 VDD.t4288 VSS 0.044149f
C18040 VDD.t2307 VSS 0.080541f
C18041 VDD.t3320 VSS 0.055186f
C18042 VDD.t2817 VSS 0.044149f
C18043 VDD.t3333 VSS 0.044149f
C18044 VDD.t2569 VSS 0.044149f
C18045 VDD.t2149 VSS 0.044149f
C18046 VDD.t2782 VSS 0.044149f
C18047 VDD.t1887 VSS 0.044149f
C18048 VDD.t2481 VSS 0.044149f
C18049 VDD.t3513 VSS 0.044149f
C18050 VDD.t2679 VSS 0.044149f
C18051 VDD.t2890 VSS 0.044149f
C18052 VDD.t1435 VSS 0.044149f
C18053 VDD.t3085 VSS 0.044149f
C18054 VDD.t3303 VSS 0.044149f
C18055 VDD.t941 VSS 0.044149f
C18056 VDD.t1020 VSS 0.033112f
C18057 VDD.n1262 VSS 0.04743f
C18058 VDD.t2755 VSS 0.055186f
C18059 VDD.t3316 VSS 0.03932f
C18060 VDD.t3230 VSS 0.026312f
C18061 VDD.t3471 VSS 0.03794f
C18062 VDD.t2946 VSS 0.040404f
C18063 VDD.t3460 VSS 0.044149f
C18064 VDD.t1160 VSS 0.022074f
C18065 VDD.t2761 VSS 0.017049f
C18066 VDD.t2763 VSS 0.036561f
C18067 VDD.t1268 VSS 0.044937f
C18068 VDD.t2750 VSS 0.041488f
C18069 VDD.t2748 VSS 0.019216f
C18070 VDD.t746 VSS 0.03252f
C18071 VDD.t1449 VSS 0.046415f
C18072 VDD.t1808 VSS 0.036659f
C18073 VDD.t3479 VSS 0.030845f
C18074 VDD.t479 VSS 0.035674f
C18075 VDD.t784 VSS 0.044149f
C18076 VDD.t778 VSS 0.020103f
C18077 VDD.t3608 VSS 0.036758f
C18078 VDD.t1151 VSS 0.03932f
C18079 VDD.n1265 VSS 0.035604f
C18080 VDD.t805 VSS 0.030845f
C18081 VDD.t1552 VSS 0.020103f
C18082 VDD.t2819 VSS 0.020103f
C18083 VDD.t759 VSS 0.02641f
C18084 VDD.t1153 VSS 0.039813f
C18085 VDD.t3624 VSS 0.020103f
C18086 VDD.t2705 VSS 0.019024f
C18087 VDD.t3620 VSS 0.030025f
C18088 VDD.t3338 VSS 0.019475f
C18089 VDD.t3622 VSS 0.025108f
C18090 VDD.t3618 VSS 0.022244f
C18091 VDD.t1779 VSS 0.033461f
C18092 VDD.t973 VSS 0.03441f
C18093 VDD.t749 VSS 0.020103f
C18094 VDD.t711 VSS 0.031141f
C18095 VDD.t2535 VSS 0.02444f
C18096 VDD.t3616 VSS 0.020103f
C18097 VDD.t3337 VSS 0.020103f
C18098 VDD.t3389 VSS 0.020103f
C18099 VDD.t2706 VSS 0.029771f
C18100 VDD.t2786 VSS 0.046707f
C18101 VDD.t1971 VSS 0.033222f
C18102 VDD.t3339 VSS 0.026544f
C18103 VDD.t279 VSS 0.027398f
C18104 VDD.t773 VSS 0.039813f
C18105 VDD.t1459 VSS 0.043557f
C18106 VDD.t3234 VSS 0.038039f
C18107 VDD.t804 VSS 0.03794f
C18108 VDD.t802 VSS 0.022938f
C18109 VDD.t34 VSS 0.028662f
C18110 VDD.t800 VSS 0.019522f
C18111 VDD.t1077 VSS 0.021436f
C18112 VDD.t811 VSS 0.037799f
C18113 VDD.t780 VSS 0.030213f
C18114 VDD.t809 VSS 0.019892f
C18115 VDD.t1068 VSS 0.020103f
C18116 VDD.t601 VSS 0.020103f
C18117 VDD.t3862 VSS 0.020103f
C18118 VDD.t3729 VSS 0.028086f
C18119 VDD.t3733 VSS 0.036265f
C18120 VDD.t2904 VSS 0.020103f
C18121 VDD.t603 VSS 0.024045f
C18122 VDD.t3393 VSS 0.022074f
C18123 VDD.t609 VSS 0.020103f
C18124 VDD.t3224 VSS 0.020103f
C18125 VDD.t3727 VSS 0.026016f
C18126 VDD.t1070 VSS 0.034294f
C18127 VDD.t4133 VSS 0.020103f
C18128 VDD.t613 VSS 0.020103f
C18129 VDD.t3024 VSS 0.034294f
C18130 VDD.t1046 VSS 0.034294f
C18131 VDD.t4145 VSS 0.024637f
C18132 VDD.t1044 VSS 0.020103f
C18133 VDD.t3388 VSS 0.02779f
C18134 VDD.t3023 VSS 0.02779f
C18135 VDD.n1272 VSS 0.023384f
C18136 VDD.n1280 VSS 0.010217f
C18137 VDD.n1281 VSS 0.015202f
C18138 VDD.n1282 VSS 0.010575f
C18139 VDD.n1285 VSS 0.017344f
C18140 VDD.n1286 VSS 0.012905f
C18141 VDD.n1291 VSS 0.014417f
C18142 VDD.n1292 VSS 0.01162f
C18143 VDD.n1298 VSS 0.01293f
C18144 VDD.n1299 VSS 0.012999f
C18145 VDD.n1300 VSS 0.011097f
C18146 VDD.n1301 VSS 0.010371f
C18147 VDD.n1304 VSS 0.019296f
C18148 VDD.n1305 VSS 0.015417f
C18149 VDD.n1312 VSS 0.01408f
C18150 VDD.n1313 VSS 0.01013f
C18151 VDD.n1329 VSS 0.01408f
C18152 VDD.n1332 VSS 0.118404f
C18153 VDD.n1333 VSS 0.017221f
C18154 VDD.n1334 VSS 0.019165f
C18155 VDD.n1335 VSS 0.019165f
C18156 VDD.n1336 VSS 0.019165f
C18157 VDD.n1337 VSS 0.019165f
C18158 VDD.n1338 VSS 0.019165f
C18159 VDD.n1339 VSS 0.127888f
C18160 VDD.t2657 VSS 0.089107f
C18161 VDD.t1502 VSS 0.088298f
C18162 VDD.t2440 VSS 0.088298f
C18163 VDD.t1158 VSS 0.088298f
C18164 VDD.t2194 VSS 0.088298f
C18165 VDD.t3037 VSS 0.088298f
C18166 VDD.t2548 VSS 0.07726f
C18167 VDD.n1340 VSS 0.04743f
C18168 VDD.t1804 VSS 0.055186f
C18169 VDD.t3068 VSS 0.088298f
C18170 VDD.t3295 VSS 0.045528f
C18171 VDD.t1330 VSS 0.025031f
C18172 VDD.t2764 VSS 0.042769f
C18173 VDD.t3911 VSS 0.059325f
C18174 VDD.t3795 VSS 0.044149f
C18175 VDD.t3293 VSS 0.021089f
C18176 VDD.t3797 VSS 0.041192f
C18177 VDD.t2262 VSS 0.027494f
C18178 VDD.t2972 VSS 0.025228f
C18179 VDD.t2384 VSS 0.022074f
C18180 VDD.t1709 VSS 0.016851f
C18181 VDD.t1711 VSS 0.019808f
C18182 VDD.t3030 VSS 0.017837f
C18183 VDD.t1939 VSS 0.034688f
C18184 VDD.t2226 VSS 0.0271f
C18185 VDD.t3546 VSS 0.023553f
C18186 VDD.t3547 VSS 0.037349f
C18187 VDD.t4135 VSS 0.03252f
C18188 VDD.t2577 VSS 0.033112f
C18189 VDD.t1029 VSS 0.040207f
C18190 VDD.t317 VSS 0.039813f
C18191 VDD.t1237 VSS 0.04001f
C18192 VDD.t1031 VSS 0.028579f
C18193 VDD.t710 VSS 0.042572f
C18194 VDD.t2438 VSS 0.047401f
C18195 VDD.t3871 VSS 0.023651f
C18196 VDD.t4165 VSS 0.03252f
C18197 VDD.t1951 VSS 0.034393f
C18198 VDD.t1950 VSS 0.024735f
C18199 VDD.t3079 VSS 0.03183f
C18200 VDD.t2410 VSS 0.036758f
C18201 VDD.t2133 VSS 0.029663f
C18202 VDD.t2131 VSS 0.028677f
C18203 VDD.t929 VSS 0.022074f
C18204 VDD.t1603 VSS 0.02444f
C18205 VDD.t137 VSS 0.051737f
C18206 VDD.t753 VSS 0.038236f
C18207 VDD.t3462 VSS 0.025425f
C18208 VDD.t1660 VSS 0.043163f
C18209 VDD.t11 VSS 0.04474f
C18210 VDD.n1346 VSS 0.050682f
C18211 VDD.n1352 VSS 0.010564f
C18212 VDD.n1353 VSS 0.01576f
C18213 VDD.n1355 VSS 0.012221f
C18214 VDD.n1356 VSS 0.018421f
C18215 VDD.n1357 VSS 0.021649f
C18216 VDD.n1360 VSS 0.015318f
C18217 VDD.n1361 VSS 0.012693f
C18218 VDD.n1362 VSS 0.011685f
C18219 VDD.n1365 VSS 0.011553f
C18220 VDD.n1367 VSS 0.013743f
C18221 VDD.n1368 VSS 0.018617f
C18222 VDD.n1369 VSS 0.01408f
C18223 VDD.n1371 VSS 0.010392f
C18224 VDD.n1372 VSS 0.118404f
C18225 VDD.n1378 VSS 0.011115f
C18226 VDD.n1379 VSS 0.010527f
C18227 VDD.n1381 VSS 0.01477f
C18228 VDD.n1382 VSS 0.012169f
C18229 VDD.n1384 VSS 0.013127f
C18230 VDD.n1385 VSS 0.113737f
C18231 VDD.t2023 VSS 0.078118f
C18232 VDD.t3400 VSS 0.044641f
C18233 VDD.t2766 VSS 0.022567f
C18234 VDD.t2650 VSS 0.03863f
C18235 VDD.t2649 VSS 0.021582f
C18236 VDD.t2442 VSS 0.044937f
C18237 VDD.t2733 VSS 0.044149f
C18238 VDD.t2170 VSS 0.016556f
C18239 VDD.t2731 VSS 0.044149f
C18240 VDD.t912 VSS 0.03252f
C18241 VDD.t2260 VSS 0.044149f
C18242 VDD.t2956 VSS 0.054496f
C18243 VDD.t2663 VSS 0.044149f
C18244 VDD.t3544 VSS 0.044149f
C18245 VDD.t3770 VSS 0.044149f
C18246 VDD.n1386 VSS 0.036885f
C18247 VDD.t2987 VSS 0.022567f
C18248 VDD.t1270 VSS 0.032619f
C18249 VDD.t3196 VSS 0.016556f
C18250 VDD.t1269 VSS 0.044641f
C18251 VDD.t2168 VSS 0.044937f
C18252 VDD.t4147 VSS 0.022074f
C18253 VDD.t2109 VSS 0.016556f
C18254 VDD.t4148 VSS 0.016556f
C18255 VDD.t2108 VSS 0.03252f
C18256 VDD.t4220 VSS 0.044937f
C18257 VDD.t1850 VSS 0.04474f
C18258 VDD.t1848 VSS 0.037349f
C18259 VDD.t2960 VSS 0.03252f
C18260 VDD.t2161 VSS 0.044149f
C18261 VDD.t3297 VSS 0.047401f
C18262 VDD.t12 VSS 0.037053f
C18263 VDD.t782 VSS 0.044149f
C18264 VDD.t738 VSS 0.048288f
C18265 VDD.t1703 VSS 0.048288f
C18266 VDD.t4131 VSS 0.023651f
C18267 VDD.t3214 VSS 0.020103f
C18268 VDD.t946 VSS 0.034491f
C18269 VDD.t2981 VSS 0.027972f
C18270 VDD.t794 VSS 0.027876f
C18271 VDD.t2983 VSS 0.019027f
C18272 VDD.t3051 VSS 0.029559f
C18273 VDD.t4014 VSS 0.030155f
C18274 VDD.t1828 VSS 0.025819f
C18275 VDD.t3283 VSS 0.02444f
C18276 VDD.t704 VSS 0.034294f
C18277 VDD.t1181 VSS 0.020103f
C18278 VDD.t1712 VSS 0.020103f
C18279 VDD.t739 VSS 0.034294f
C18280 VDD.t1826 VSS 0.02444f
C18281 VDD.t3281 VSS 0.025819f
C18282 VDD.t3216 VSS 0.034118f
C18283 VDD.t2223 VSS 0.030017f
C18284 VDD.t945 VSS 0.019475f
C18285 VDD.t2671 VSS 0.019475f
C18286 VDD.t2225 VSS 0.02253f
C18287 VDD.t906 VSS 0.018927f
C18288 VDD.t2397 VSS 0.034572f
C18289 VDD.t713 VSS 0.025228f
C18290 VDD.t1941 VSS 0.02641f
C18291 VDD.t3287 VSS 0.028776f
C18292 VDD.t3218 VSS 0.021089f
C18293 VDD.t3285 VSS 0.020103f
C18294 VDD.t948 VSS 0.023848f
C18295 VDD.t3217 VSS 0.040207f
C18296 VDD.t2470 VSS 0.038433f
C18297 VDD.n1393 VSS 0.037575f
C18298 VDD.n1400 VSS 0.016303f
C18299 VDD.n1401 VSS 0.013941f
C18300 VDD.n1404 VSS 0.01515f
C18301 VDD.n1405 VSS 0.010295f
C18302 VDD.n1406 VSS 0.012711f
C18303 VDD.n1408 VSS 0.02025f
C18304 VDD.n1409 VSS 0.024323f
C18305 VDD.n1411 VSS 0.014181f
C18306 VDD.n1412 VSS 0.014684f
C18307 VDD.n1413 VSS 0.013884f
C18308 VDD.n1414 VSS 0.014181f
C18309 VDD.n1416 VSS 0.011903f
C18310 VDD.n1417 VSS 0.01094f
C18311 VDD.n1418 VSS 0.118404f
C18312 VDD.n1419 VSS 0.378819f
C18313 VDD.n1420 VSS 0.010228f
C18314 VDD.n1425 VSS 0.012807f
C18315 VDD.n1427 VSS 0.012511f
C18316 VDD.n1428 VSS 0.012417f
C18317 VDD.n1433 VSS 0.012361f
C18318 VDD.n1439 VSS 0.012369f
C18319 VDD.n1442 VSS 0.012916f
C18320 VDD.n1457 VSS 0.011924f
C18321 VDD.n1460 VSS 0.012711f
C18322 VDD.n1462 VSS 0.012257f
C18323 VDD.n1463 VSS 0.011074f
C18324 VDD.n1467 VSS 0.012527f
C18325 VDD.n1468 VSS 0.010296f
C18326 VDD.n1474 VSS 0.013806f
C18327 VDD.n1476 VSS 0.011383f
C18328 VDD.n1481 VSS 0.013031f
C18329 VDD.n1482 VSS 0.231769f
C18330 VDD.n1483 VSS 0.010392f
C18331 VDD.n1488 VSS 0.010337f
C18332 VDD.n1489 VSS 0.010828f
C18333 VDD.n1493 VSS 0.010417f
C18334 VDD.n1494 VSS 0.011383f
C18335 VDD.n1498 VSS 0.01723f
C18336 VDD.n1499 VSS 0.02136f
C18337 VDD.n1501 VSS 0.014613f
C18338 VDD.n1502 VSS 0.01603f
C18339 VDD.n1504 VSS 0.011429f
C18340 VDD.n1505 VSS 0.015065f
C18341 VDD.n1507 VSS 0.011999f
C18342 VDD.n1508 VSS 0.036984f
C18343 VDD.t3628 VSS 0.028184f
C18344 VDD.t2332 VSS 0.02444f
C18345 VDD.t2184 VSS 0.022074f
C18346 VDD.t2334 VSS 0.025228f
C18347 VDD.t2349 VSS 0.044149f
C18348 VDD.t2347 VSS 0.044149f
C18349 VDD.t2343 VSS 0.044149f
C18350 VDD.t2345 VSS 0.044149f
C18351 VDD.t2340 VSS 0.044149f
C18352 VDD.t457 VSS 0.044149f
C18353 VDD.t459 VSS 0.044149f
C18354 VDD.t451 VSS 0.044149f
C18355 VDD.t453 VSS 0.044149f
C18356 VDD.t455 VSS 0.044149f
C18357 VDD.t619 VSS 0.044149f
C18358 VDD.t447 VSS 0.028381f
C18359 VDD.t2293 VSS 0.022074f
C18360 VDD.t449 VSS 0.023651f
C18361 VDD.t3768 VSS 0.038942f
C18362 VDD.n1509 VSS 0.105436f
C18363 VDD.n1524 VSS 0.429013f
C18364 VDD.n1525 VSS 0.118404f
C18365 VDD.n1528 VSS 0.010053f
C18366 VDD.n1529 VSS 0.017433f
C18367 VDD.n1535 VSS 0.010055f
C18368 VDD.n1536 VSS 0.014602f
C18369 VDD.n1538 VSS 0.010013f
C18370 VDD.n1540 VSS 0.013771f
C18371 VDD.n1541 VSS 0.014702f
C18372 VDD.n1545 VSS 0.021224f
C18373 VDD.n1546 VSS 0.021887f
C18374 VDD.n1547 VSS 0.013028f
C18375 VDD.n1548 VSS 0.010261f
C18376 VDD.n1549 VSS 0.011222f
C18377 VDD.n1554 VSS 0.013194f
C18378 VDD.n1555 VSS 0.010721f
C18379 VDD.n1557 VSS 0.020143f
C18380 VDD.n1558 VSS 0.011266f
C18381 VDD.n1559 VSS 0.011803f
C18382 VDD.n1560 VSS 0.010982f
C18383 VDD.n1562 VSS 0.014274f
C18384 VDD.n1565 VSS 0.017453f
C18385 VDD.n1566 VSS 0.01939f
C18386 VDD.n1568 VSS 0.011876f
C18387 VDD.n1569 VSS 0.011549f
C18388 VDD.n1570 VSS 0.013725f
C18389 VDD.n1575 VSS 0.118404f
C18390 VDD.n1576 VSS 0.118404f
C18391 VDD.n1577 VSS 0.014061f
C18392 VDD.n1578 VSS 0.017764f
C18393 VDD.n1579 VSS 0.010888f
C18394 VDD.n1580 VSS 0.014162f
C18395 VDD.n1581 VSS 0.014741f
C18396 VDD.n1582 VSS 0.017471f
C18397 VDD.n1583 VSS 0.011002f
C18398 VDD.n1584 VSS 0.014118f
C18399 VDD.n1585 VSS 0.014246f
C18400 VDD.n1586 VSS 0.010571f
C18401 VDD.n1587 VSS 0.014892f
C18402 VDD.n1591 VSS 0.012579f
C18403 VDD.n1593 VSS 0.010742f
C18404 VDD.n1596 VSS 0.014778f
C18405 VDD.n1597 VSS 0.039053f
C18406 VDD.t3017 VSS 0.030155f
C18407 VDD.t3511 VSS 0.033604f
C18408 VDD.t876 VSS 0.022764f
C18409 VDD.t2353 VSS 0.020793f
C18410 VDD.t509 VSS 0.021385f
C18411 VDD.t442 VSS 0.021385f
C18412 VDD.t2052 VSS 0.023158f
C18413 VDD.t3019 VSS 0.023158f
C18414 VDD.t943 VSS 0.047302f
C18415 VDD.t1101 VSS 0.028671f
C18416 VDD.t2745 VSS 0.022912f
C18417 VDD.t1513 VSS 0.027876f
C18418 VDD.t3652 VSS 0.035306f
C18419 VDD.t1495 VSS 0.034391f
C18420 VDD.t531 VSS 0.025622f
C18421 VDD.t3507 VSS 0.031141f
C18422 VDD.t1928 VSS 0.022074f
C18423 VDD.t3509 VSS 0.020103f
C18424 VDD.t2742 VSS 0.02917f
C18425 VDD.t944 VSS 0.035772f
C18426 VDD.t2328 VSS 0.020103f
C18427 VDD.t4028 VSS 0.03252f
C18428 VDD.t1483 VSS 0.034294f
C18429 VDD.t2743 VSS 0.016556f
C18430 VDD.t1485 VSS 0.020103f
C18431 VDD.t360 VSS 0.039911f
C18432 VDD.n1598 VSS 0.038462f
C18433 VDD.t3782 VSS 0.021582f
C18434 VDD.t3780 VSS 0.02099f
C18435 VDD.t783 VSS 0.022074f
C18436 VDD.t3766 VSS 0.055186f
C18437 VDD.t529 VSS 0.088101f
C18438 VDD.t2117 VSS 0.057354f
C18439 VDD.t792 VSS 0.02986f
C18440 VDD.t1081 VSS 0.025721f
C18441 VDD.t3114 VSS 0.019216f
C18442 VDD.t3116 VSS 0.04474f
C18443 VDD.t2389 VSS 0.044937f
C18444 VDD.t3189 VSS 0.03252f
C18445 VDD.t2508 VSS 0.016556f
C18446 VDD.t3190 VSS 0.016556f
C18447 VDD.t2507 VSS 0.022074f
C18448 VDD.t155 VSS 0.044937f
C18449 VDD.t1927 VSS 0.047598f
C18450 VDD.t3429 VSS 0.016556f
C18451 VDD.t1925 VSS 0.024045f
C18452 VDD.t1074 VSS 0.022074f
C18453 VDD.t2408 VSS 0.020103f
C18454 VDD.t796 VSS 0.044641f
C18455 VDD.n1604 VSS 0.052061f
C18456 VDD.t3542 VSS 0.033112f
C18457 VDD.t2930 VSS 0.034294f
C18458 VDD.t1973 VSS 0.022074f
C18459 VDD.t4222 VSS 0.018822f
C18460 VDD.t4224 VSS 0.017837f
C18461 VDD.t515 VSS 0.025721f
C18462 VDD.t3540 VSS 0.041685f
C18463 VDD.t2198 VSS 0.020103f
C18464 VDD.t3362 VSS 0.015671f
C18465 VDD.t2199 VSS 0.029882f
C18466 VDD.t3357 VSS 0.027113f
C18467 VDD.t1956 VSS 0.027685f
C18468 VDD.t1958 VSS 0.016229f
C18469 VDD.t2932 VSS 0.033724f
C18470 VDD.t467 VSS 0.042902f
C18471 VDD.t4035 VSS 0.025031f
C18472 VDD.t4036 VSS 0.022666f
C18473 VDD.t2892 VSS 0.026213f
C18474 VDD.t3360 VSS 0.02641f
C18475 VDD.t2788 VSS 0.020103f
C18476 VDD.t3361 VSS 0.0339f
C18477 VDD.t3710 VSS 0.028776f
C18478 VDD.t3834 VSS 0.032323f
C18479 VDD.t1107 VSS 0.025622f
C18480 VDD.t3358 VSS 0.022074f
C18481 VDD.t358 VSS 0.051188f
C18482 VDD.n1612 VSS 0.109173f
C18483 VDD.n1614 VSS 0.013963f
C18484 VDD.n1615 VSS 0.013137f
C18485 VDD.n1616 VSS 0.010165f
C18486 VDD.n1617 VSS 0.014188f
C18487 VDD.n1618 VSS 0.015335f
C18488 VDD.n1619 VSS 0.012139f
C18489 VDD.n1624 VSS 0.014586f
C18490 VDD.n1626 VSS 0.010092f
C18491 VDD.n1627 VSS 0.012906f
C18492 VDD.n1628 VSS 0.010818f
C18493 VDD.n1629 VSS 0.015272f
C18494 VDD.n1630 VSS 0.015669f
C18495 VDD.n1631 VSS 0.020132f
C18496 VDD.n1632 VSS 0.018879f
C18497 VDD.n1633 VSS 0.018199f
C18498 VDD.n1634 VSS 0.011538f
C18499 VDD.n1636 VSS 0.010993f
C18500 VDD.n1637 VSS 0.013701f
C18501 VDD.n1642 VSS 0.118404f
C18502 VDD.n1643 VSS 0.118404f
C18503 VDD.n1653 VSS 0.014583f
C18504 VDD.n1654 VSS 0.013217f
C18505 VDD.n1656 VSS 0.012939f
C18506 VDD.n1657 VSS 0.014631f
C18507 VDD.n1660 VSS 0.014211f
C18508 VDD.n1661 VSS 0.013507f
C18509 VDD.n1662 VSS 0.012956f
C18510 VDD.n1663 VSS 0.012173f
C18511 VDD.n1664 VSS 0.012036f
C18512 VDD.n1665 VSS 0.011689f
C18513 VDD.n1668 VSS 0.013532f
C18514 VDD.n1669 VSS 0.036582f
C18515 VDD.t537 VSS 0.029104f
C18516 VDD.t2687 VSS 0.038932f
C18517 VDD.t28 VSS 0.02641f
C18518 VDD.t3840 VSS 0.020103f
C18519 VDD.t3222 VSS 0.034294f
C18520 VDD.t2689 VSS 0.036955f
C18521 VDD.t2918 VSS 0.038532f
C18522 VDD.t2916 VSS 0.023355f
C18523 VDD.t2406 VSS 0.021385f
C18524 VDD.t3819 VSS 0.020793f
C18525 VDD.t2920 VSS 0.020103f
C18526 VDD.t1702 VSS 0.022074f
C18527 VDD.t2914 VSS 0.020103f
C18528 VDD.t1869 VSS 0.022074f
C18529 VDD.t575 VSS 0.026706f
C18530 VDD.t856 VSS 0.033112f
C18531 VDD.t3590 VSS 0.022074f
C18532 VDD.t854 VSS 0.020103f
C18533 VDD.t3866 VSS 0.022074f
C18534 VDD.t573 VSS 0.02444f
C18535 VDD.t1109 VSS 0.022074f
C18536 VDD.t571 VSS 0.032717f
C18537 VDD.t850 VSS 0.039419f
C18538 VDD.t3993 VSS 0.022074f
C18539 VDD.t852 VSS 0.023651f
C18540 VDD.t1263 VSS 0.022074f
C18541 VDD.t858 VSS 0.042033f
C18542 VDD.n1670 VSS 0.114915f
C18543 VDD.n1675 VSS 0.013457f
C18544 VDD.n1676 VSS 0.014154f
C18545 VDD.n1679 VSS 0.011444f
C18546 VDD.n1683 VSS 0.118404f
C18547 VDD.n1684 VSS 0.118404f
C18548 VDD.n1689 VSS 0.016365f
C18549 VDD.n1691 VSS 0.014938f
C18550 VDD.n1692 VSS 0.014999f
C18551 VDD.n1693 VSS 0.015772f
C18552 VDD.n1694 VSS 0.016308f
C18553 VDD.n1695 VSS 0.010468f
C18554 VDD.n1696 VSS 0.011021f
C18555 VDD.n1698 VSS 0.011151f
C18556 VDD.n1699 VSS 0.013532f
C18557 VDD.n1712 VSS 0.010077f
C18558 VDD.n1715 VSS 0.010903f
C18559 VDD.n1718 VSS 0.015886f
C18560 VDD.n1724 VSS 0.014264f
C18561 VDD.n1725 VSS 0.010322f
C18562 VDD.n1729 VSS 0.010371f
C18563 VDD.n1735 VSS 0.01408f
C18564 VDD.n1740 VSS 0.010392f
C18565 VDD.n1741 VSS 0.118404f
C18566 VDD.n1742 VSS 0.118404f
C18567 VDD.n1748 VSS 0.014846f
C18568 VDD.n1773 VSS 0.01065f
C18569 VDD.n1774 VSS 0.013806f
C18570 VDD.n1775 VSS 0.025355f
C18571 VDD.t599 VSS 0.039221f
C18572 VDD.t607 VSS 0.035083f
C18573 VDD.t275 VSS 0.033112f
C18574 VDD.t1966 VSS 0.031141f
C18575 VDD.t139 VSS 0.034294f
C18576 VDD.t1798 VSS 0.024045f
C18577 VDD.t141 VSS 0.020103f
C18578 VDD.t1806 VSS 0.020103f
C18579 VDD.t151 VSS 0.020103f
C18580 VDD.t1968 VSS 0.024045f
C18581 VDD.t143 VSS 0.020103f
C18582 VDD.t2121 VSS 0.023651f
C18583 VDD.t689 VSS 0.031141f
C18584 VDD.t481 VSS 0.024045f
C18585 VDD.t699 VSS 0.021286f
C18586 VDD.t687 VSS 0.033787f
C18587 VDD.t1477 VSS 0.022397f
C18588 VDD.t697 VSS 0.027876f
C18589 VDD.t1965 VSS 0.019475f
C18590 VDD.t661 VSS 0.025501f
C18591 VDD.t695 VSS 0.027116f
C18592 VDD.t1807 VSS 0.020103f
C18593 VDD.t659 VSS 0.020103f
C18594 VDD.t3959 VSS 0.024045f
C18595 VDD.t663 VSS 0.02444f
C18596 VDD.t523 VSS 0.02375f
C18597 VDD.t2906 VSS 0.050949f
C18598 VDD.n1776 VSS 0.037575f
C18599 VDD.t3961 VSS 0.028184f
C18600 VDD.t43 VSS 0.035772f
C18601 VDD.t125 VSS 0.024045f
C18602 VDD.t117 VSS 0.024045f
C18603 VDD.t119 VSS 0.020103f
C18604 VDD.t41 VSS 0.020103f
C18605 VDD.t621 VSS 0.024045f
C18606 VDD.t121 VSS 0.024045f
C18607 VDD.t123 VSS 0.023651f
C18608 VDD.t352 VSS 0.023651f
C18609 VDD.t2608 VSS 0.024045f
C18610 VDD.t319 VSS 0.024045f
C18611 VDD.t2610 VSS 0.020103f
C18612 VDD.t388 VSS 0.020103f
C18613 VDD.t2634 VSS 0.024045f
C18614 VDD.t354 VSS 0.024045f
C18615 VDD.t2606 VSS 0.020103f
C18616 VDD.t386 VSS 0.020103f
C18617 VDD.t2614 VSS 0.024045f
C18618 VDD.t347 VSS 0.024045f
C18619 VDD.t2638 VSS 0.020103f
C18620 VDD.t321 VSS 0.020103f
C18621 VDD.t2612 VSS 0.024045f
C18622 VDD.t390 VSS 0.024045f
C18623 VDD.t2636 VSS 0.048091f
C18624 VDD.t4118 VSS 0.044937f
C18625 VDD.t3299 VSS 0.02444f
C18626 VDD.t638 VSS 0.023651f
C18627 VDD.t1222 VSS 0.020103f
C18628 VDD.t1891 VSS 0.030155f
C18629 VDD.n1788 VSS 0.039053f
C18630 VDD.t2952 VSS 0.033604f
C18631 VDD.t2019 VSS 0.034294f
C18632 VDD.t3039 VSS 0.022074f
C18633 VDD.t2566 VSS 0.019315f
C18634 VDD.t2568 VSS 0.017344f
C18635 VDD.t520 VSS 0.025228f
C18636 VDD.t2950 VSS 0.044149f
C18637 VDD.t920 VSS 0.020103f
C18638 VDD.t3073 VSS 0.016616f
C18639 VDD.t921 VSS 0.02886f
C18640 VDD.t3493 VSS 0.031504f
C18641 VDD.t1830 VSS 0.027876f
C18642 VDD.t1025 VSS 0.039458f
C18643 VDD.t3242 VSS 0.034405f
C18644 VDD.t475 VSS 0.023651f
C18645 VDD.t4022 VSS 0.031141f
C18646 VDD.t2999 VSS 0.031141f
C18647 VDD.t3496 VSS 0.040207f
C18648 VDD.t3072 VSS 0.040207f
C18649 VDD.t1525 VSS 0.032323f
C18650 VDD.t4065 VSS 0.034294f
C18651 VDD.t3494 VSS 0.042178f
C18652 VDD.t364 VSS 0.051145f
C18653 VDD.n1795 VSS 0.104437f
C18654 VDD.n1797 VSS 0.019575f
C18655 VDD.n1798 VSS 0.01512f
C18656 VDD.n1800 VSS 0.012422f
C18657 VDD.n1801 VSS 0.015669f
C18658 VDD.n1802 VSS 0.012481f
C18659 VDD.n1807 VSS 0.017515f
C18660 VDD.n1808 VSS 0.011818f
C18661 VDD.n1824 VSS 0.011383f
C18662 VDD.n1829 VSS 0.011151f
C18663 VDD.n1830 VSS 0.01163f
C18664 VDD.n1835 VSS 0.010885f
C18665 VDD.n1836 VSS 0.118404f
C18666 VDD.n1837 VSS 0.118404f
C18667 VDD.n1840 VSS 0.013247f
C18668 VDD.n1842 VSS 0.012859f
C18669 VDD.n1843 VSS 0.013643f
C18670 VDD.n1845 VSS 0.020759f
C18671 VDD.n1846 VSS 0.012465f
C18672 VDD.n1847 VSS 0.015007f
C18673 VDD.n1848 VSS 0.0184f
C18674 VDD.n1849 VSS 0.015272f
C18675 VDD.n1850 VSS 0.015272f
C18676 VDD.n1851 VSS 0.020303f
C18677 VDD.n1852 VSS 0.016928f
C18678 VDD.n1856 VSS 0.013532f
C18679 VDD.n1857 VSS 0.037575f
C18680 VDD.t2382 VSS 0.028874f
C18681 VDD.t499 VSS 0.021385f
C18682 VDD.t844 VSS 0.02444f
C18683 VDD.t3194 VSS 0.02444f
C18684 VDD.t1257 VSS 0.020103f
C18685 VDD.t4044 VSS 0.048334f
C18686 VDD.t1489 VSS 0.03094f
C18687 VDD.t1175 VSS 0.023676f
C18688 VDD.t1177 VSS 0.025585f
C18689 VDD.t1493 VSS 0.021353f
C18690 VDD.t1173 VSS 0.034252f
C18691 VDD.t477 VSS 0.022074f
C18692 VDD.t1171 VSS 0.027593f
C18693 VDD.t83 VSS 0.025622f
C18694 VDD.t2136 VSS 0.022074f
C18695 VDD.t67 VSS 0.020103f
C18696 VDD.t1492 VSS 0.02168f
C18697 VDD.t4045 VSS 0.020498f
C18698 VDD.t85 VSS 0.020103f
C18699 VDD.t910 VSS 0.022074f
C18700 VDD.t69 VSS 0.02444f
C18701 VDD.t71 VSS 0.031929f
C18702 VDD.t1490 VSS 0.022074f
C18703 VDD.t416 VSS 0.020103f
C18704 VDD.t2626 VSS 0.022074f
C18705 VDD.t65 VSS 0.036265f
C18706 VDD.t63 VSS 0.031929f
C18707 VDD.t4274 VSS 0.038942f
C18708 VDD.n1858 VSS 0.100569f
C18709 VDD.n1859 VSS 0.0108f
C18710 VDD.n1864 VSS 0.012965f
C18711 VDD.n1869 VSS 0.013784f
C18712 VDD.n1870 VSS 0.011323f
C18713 VDD.n1871 VSS 0.118404f
C18714 VDD.n1872 VSS 0.118404f
C18715 VDD.n1877 VSS 0.06795f
C18716 VDD.n1879 VSS 0.016867f
C18717 VDD.n1880 VSS 0.014999f
C18718 VDD.n1881 VSS 0.014938f
C18719 VDD.n1882 VSS 0.015485f
C18720 VDD.n1885 VSS 0.014724f
C18721 VDD.n1886 VSS 0.021416f
C18722 VDD.n1888 VSS 0.010157f
C18723 VDD.n1891 VSS 0.010108f
C18724 VDD.n1894 VSS 0.012063f
C18725 VDD.n1897 VSS 0.011565f
C18726 VDD.n1898 VSS 0.013665f
C18727 VDD.n1899 VSS 0.014897f
C18728 VDD.n1900 VSS 0.017118f
C18729 VDD.n1902 VSS 0.012072f
C18730 VDD.n1904 VSS 0.011312f
C18731 VDD.n1905 VSS 0.014556f
C18732 VDD.n1906 VSS 0.012577f
C18733 VDD.n1908 VSS 0.011001f
C18734 VDD.n1909 VSS 0.011015f
C18735 VDD.n1910 VSS 0.011015f
C18736 VDD.n1911 VSS 0.01508f
C18737 VDD.n1912 VSS 0.013647f
C18738 VDD.n1913 VSS 0.01408f
C18739 VDD.n1914 VSS 0.01013f
C18740 VDD.n1920 VSS 0.118404f
C18741 VDD.n1921 VSS 0.118404f
C18742 VDD.n1927 VSS 0.01013f
C18743 VDD.n1928 VSS 0.01408f
C18744 VDD.n1929 VSS 0.013647f
C18745 VDD.n1930 VSS 0.01508f
C18746 VDD.n1931 VSS 0.014669f
C18747 VDD.n1932 VSS 0.011236f
C18748 VDD.n1933 VSS 0.010381f
C18749 VDD.n1937 VSS 0.011057f
C18750 VDD.n1938 VSS 0.015575f
C18751 VDD.n1939 VSS 0.01233f
C18752 VDD.n1943 VSS 0.010446f
C18753 VDD.n1945 VSS 0.010742f
C18754 VDD.n1948 VSS 0.013642f
C18755 VDD.n1949 VSS 0.037611f
C18756 VDD.t723 VSS 0.029663f
C18757 VDD.t4009 VSS 0.031141f
C18758 VDD.t2080 VSS 0.03321f
C18759 VDD.t1279 VSS 0.021188f
C18760 VDD.t3047 VSS 0.020103f
C18761 VDD.t3750 VSS 0.020103f
C18762 VDD.t539 VSS 0.020103f
C18763 VDD.t2866 VSS 0.02444f
C18764 VDD.t4007 VSS 0.025524f
C18765 VDD.t3582 VSS 0.028874f
C18766 VDD.t1276 VSS 0.029303f
C18767 VDD.t277 VSS 0.019323f
C18768 VDD.t3473 VSS 0.02864f
C18769 VDD.t4030 VSS 0.042336f
C18770 VDD.t441 VSS 0.034186f
C18771 VDD.t492 VSS 0.020103f
C18772 VDD.t412 VSS 0.020892f
C18773 VDD.t1203 VSS 0.030352f
C18774 VDD.t1463 VSS 0.027593f
C18775 VDD.t410 VSS 0.020103f
C18776 VDD.t3474 VSS 0.020103f
C18777 VDD.t439 VSS 0.020103f
C18778 VDD.t3583 VSS 0.022863f
C18779 VDD.t2948 VSS 0.039024f
C18780 VDD.t1963 VSS 0.034294f
C18781 VDD.t3475 VSS 0.02444f
C18782 VDD.t3983 VSS 0.020103f
C18783 VDD.t2618 VSS 0.030155f
C18784 VDD.n1950 VSS 0.039546f
C18785 VDD.t788 VSS 0.029465f
C18786 VDD.t2311 VSS 0.032422f
C18787 VDD.t2562 VSS 0.029663f
C18788 VDD.t351 VSS 0.020103f
C18789 VDD.t787 VSS 0.030648f
C18790 VDD.t1092 VSS 0.051047f
C18791 VDD.t3595 VSS 0.043163f
C18792 VDD.t2097 VSS 0.03252f
C18793 VDD.t3570 VSS 0.022074f
C18794 VDD.t1735 VSS 0.016556f
C18795 VDD.t3569 VSS 0.016556f
C18796 VDD.t1734 VSS 0.044937f
C18797 VDD.t1947 VSS 0.044937f
C18798 VDD.t1543 VSS 0.016556f
C18799 VDD.t1948 VSS 0.016556f
C18800 VDD.t1541 VSS 0.022074f
C18801 VDD.t1403 VSS 0.03252f
C18802 VDD.t2436 VSS 0.040995f
C18803 VDD.t963 VSS 0.048879f
C18804 VDD.t3815 VSS 0.040207f
C18805 VDD.t1773 VSS 0.020596f
C18806 VDD.t485 VSS 0.020103f
C18807 VDD.t1836 VSS 0.02917f
C18808 VDD.t2142 VSS 0.031633f
C18809 VDD.n1957 VSS 0.043981f
C18810 VDD.t992 VSS 0.030155f
C18811 VDD.t1287 VSS 0.034294f
C18812 VDD.t1935 VSS 0.023651f
C18813 VDD.t2376 VSS 0.020103f
C18814 VDD.t501 VSS 0.043656f
C18815 VDD.t994 VSS 0.032422f
C18816 VDD.t1664 VSS 0.020103f
C18817 VDD.t1880 VSS 0.022074f
C18818 VDD.t1670 VSS 0.029602f
C18819 VDD.t3363 VSS 0.020896f
C18820 VDD.t1668 VSS 0.023676f
C18821 VDD.t1666 VSS 0.025585f
C18822 VDD.t1093 VSS 0.021353f
C18823 VDD.t313 VSS 0.034252f
C18824 VDD.t517 VSS 0.022074f
C18825 VDD.t309 VSS 0.027593f
C18826 VDD.t303 VSS 0.025622f
C18827 VDD.t1120 VSS 0.022074f
C18828 VDD.t301 VSS 0.020103f
C18829 VDD.t3366 VSS 0.02168f
C18830 VDD.t1879 VSS 0.020498f
C18831 VDD.t307 VSS 0.020103f
C18832 VDD.t2176 VSS 0.022074f
C18833 VDD.t315 VSS 0.02444f
C18834 VDD.t311 VSS 0.031929f
C18835 VDD.t3364 VSS 0.022074f
C18836 VDD.t305 VSS 0.020103f
C18837 VDD.t2630 VSS 0.038942f
C18838 VDD.n1967 VSS 0.105436f
C18839 VDD.n1971 VSS 0.012965f
C18840 VDD.n1976 VSS 0.013184f
C18841 VDD.n1977 VSS 0.010869f
C18842 VDD.n1983 VSS 0.017077f
C18843 VDD.n1984 VSS 0.014825f
C18844 VDD.n1985 VSS 0.015907f
C18845 VDD.n1987 VSS 0.015272f
C18846 VDD.n1988 VSS 0.015272f
C18847 VDD.n1989 VSS 0.01543f
C18848 VDD.n1990 VSS 0.020068f
C18849 VDD.n1992 VSS 0.012984f
C18850 VDD.n1995 VSS 0.015469f
C18851 VDD.n1996 VSS 0.014263f
C18852 VDD.n1998 VSS 0.012545f
C18853 VDD.n1999 VSS 0.011159f
C18854 VDD.n2000 VSS 0.118404f
C18855 VDD.n2001 VSS 0.118404f
C18856 VDD.n2003 VSS 0.013101f
C18857 VDD.n2004 VSS 0.020409f
C18858 VDD.n2005 VSS 0.015549f
C18859 VDD.n2008 VSS 0.019718f
C18860 VDD.n2009 VSS 0.014408f
C18861 VDD.n2010 VSS 0.016912f
C18862 VDD.n2011 VSS 0.015669f
C18863 VDD.n2012 VSS 0.012084f
C18864 VDD.n2013 VSS 0.010742f
C18865 VDD.n2017 VSS 0.012612f
C18866 VDD.n2018 VSS 0.013123f
C18867 VDD.n2023 VSS 0.037575f
C18868 VDD.t2924 VSS 0.033604f
C18869 VDD.t1867 VSS 0.020103f
C18870 VDD.t486 VSS 0.022074f
C18871 VDD.t2588 VSS 0.02444f
C18872 VDD.t3690 VSS 0.016556f
C18873 VDD.t2587 VSS 0.020103f
C18874 VDD.t1 VSS 0.041731f
C18875 VDD.t2188 VSS 0.031608f
C18876 VDD.t1192 VSS 0.018998f
C18877 VDD.t1193 VSS 0.024917f
C18878 VDD.t2241 VSS 0.031561f
C18879 VDD.t3232 VSS 0.034339f
C18880 VDD.t461 VSS 0.042079f
C18881 VDD.t2556 VSS 0.036462f
C18882 VDD.t644 VSS 0.020103f
C18883 VDD.t2191 VSS 0.034885f
C18884 VDD.t0 VSS 0.029367f
C18885 VDD.t4063 VSS 0.020103f
C18886 VDD.t1548 VSS 0.045134f
C18887 VDD.t2189 VSS 0.037448f
C18888 VDD.t4205 VSS 0.020103f
C18889 VDD.t2616 VSS 0.020103f
C18890 VDD.t3486 VSS 0.027199f
C18891 VDD.t3638 VSS 0.060964f
C18892 VDD.n2024 VSS 0.114603f
C18893 VDD.n2025 VSS 0.011361f
C18894 VDD.n2027 VSS 0.017084f
C18895 VDD.n2028 VSS 0.01939f
C18896 VDD.n2030 VSS 0.013986f
C18897 VDD.n2031 VSS 0.017291f
C18898 VDD.n2032 VSS 0.118404f
C18899 VDD.n2033 VSS 0.118404f
C18900 VDD.n2038 VSS 0.016119f
C18901 VDD.n2040 VSS 0.010092f
C18902 VDD.n2041 VSS 0.014029f
C18903 VDD.n2042 VSS 0.010211f
C18904 VDD.n2044 VSS 0.017494f
C18905 VDD.n2045 VSS 0.013137f
C18906 VDD.n2047 VSS 0.011546f
C18907 VDD.n2048 VSS 0.010659f
C18908 VDD.n2049 VSS 0.011769f
C18909 VDD.n2050 VSS 0.013094f
C18910 VDD.n2052 VSS 0.010742f
C18911 VDD.n2054 VSS 0.010692f
C18912 VDD.n2055 VSS 0.013287f
C18913 VDD.n2056 VSS 0.010742f
C18914 VDD.n2057 VSS 0.010702f
C18915 VDD.n2058 VSS 0.011077f
C18916 VDD.n2059 VSS 0.011686f
C18917 VDD.n2060 VSS 0.015461f
C18918 VDD.n2063 VSS 0.018993f
C18919 VDD.n2067 VSS 0.012648f
C18920 VDD.n2068 VSS 0.015714f
C18921 VDD.n2069 VSS 0.019165f
C18922 VDD.n2070 VSS 0.019165f
C18923 VDD.n2071 VSS 0.019165f
C18924 VDD.n2072 VSS 0.019165f
C18925 VDD.n2073 VSS 0.017084f
C18926 VDD.n2074 VSS 0.01408f
C18927 VDD.n2075 VSS 0.01013f
C18928 VDD.n2081 VSS 0.118404f
C18929 VDD.n2082 VSS 0.118404f
C18930 VDD.n2088 VSS 0.01013f
C18931 VDD.n2089 VSS 0.01408f
C18932 VDD.n2090 VSS 0.017084f
C18933 VDD.n2091 VSS 0.019165f
C18934 VDD.n2092 VSS 0.019165f
C18935 VDD.n2093 VSS 0.019165f
C18936 VDD.n2094 VSS 0.019165f
C18937 VDD.n2095 VSS 0.019165f
C18938 VDD.n2096 VSS 0.019165f
C18939 VDD.n2097 VSS 0.019165f
C18940 VDD.n2098 VSS 0.01013f
C18941 VDD.n2100 VSS 0.016392f
C18942 VDD.n2101 VSS 0.015274f
C18943 VDD.n2102 VSS 0.014682f
C18944 VDD.n2103 VSS 0.04743f
C18945 VDD.t2719 VSS 0.040207f
C18946 VDD.t718 VSS 0.043557f
C18947 VDD.t2282 VSS 0.038433f
C18948 VDD.t2285 VSS 0.044149f
C18949 VDD.t1648 VSS 0.044149f
C18950 VDD.t1646 VSS 0.044149f
C18951 VDD.t1638 VSS 0.044149f
C18952 VDD.t1650 VSS 0.044149f
C18953 VDD.t1642 VSS 0.044149f
C18954 VDD.t1636 VSS 0.044149f
C18955 VDD.t1640 VSS 0.023651f
C18956 VDD.t2737 VSS 0.024045f
C18957 VDD.t1644 VSS 0.024045f
C18958 VDD.t2734 VSS 0.023651f
C18959 VDD.t761 VSS 0.044149f
C18960 VDD.t715 VSS 0.044149f
C18961 VDD.t771 VSS 0.034393f
C18962 VDD.t15 VSS 0.024045f
C18963 VDD.t719 VSS 0.020103f
C18964 VDD.t3598 VSS 0.039221f
C18965 VDD.n2104 VSS 0.049302f
C18966 VDD.n2109 VSS 0.023124f
C18967 VDD.t937 VSS 0.041028f
C18968 VDD.t3125 VSS 0.042769f
C18969 VDD.t4193 VSS 0.031535f
C18970 VDD.t3123 VSS 0.022074f
C18971 VDD.t4195 VSS 0.02444f
C18972 VDD.t648 VSS 0.028381f
C18973 VDD.t2257 VSS 0.037743f
C18974 VDD.t2428 VSS 0.039714f
C18975 VDD.t3501 VSS 0.024538f
C18976 VDD.t3588 VSS 0.016556f
C18977 VDD.t3503 VSS 0.024045f
C18978 VDD.t3490 VSS 0.030057f
C18979 VDD.t3273 VSS 0.034984f
C18980 VDD.t1883 VSS 0.031436f
C18981 VDD.t1881 VSS 0.021483f
C18982 VDD.t4107 VSS 0.025031f
C18983 VDD.t2238 VSS 0.027593f
C18984 VDD.t2244 VSS 0.036462f
C18985 VDD.t2825 VSS 0.058438f
C18986 VDD.t503 VSS 0.034294f
C18987 VDD.t1908 VSS 0.024932f
C18988 VDD.t488 VSS 0.03932f
C18989 VDD.t536 VSS 0.02444f
C18990 VDD.t2827 VSS 0.025326f
C18991 VDD.t1454 VSS 0.031141f
C18992 VDD.n2114 VSS 0.032969f
C18993 VDD.t1676 VSS 0.033123f
C18994 VDD.t507 VSS 0.041784f
C18995 VDD.t2426 VSS 0.031141f
C18996 VDD.t2434 VSS 0.023651f
C18997 VDD.t3714 VSS 0.020103f
C18998 VDD.t2035 VSS 0.02917f
C18999 VDD.t1453 VSS 0.029367f
C19000 VDD.t471 VSS 0.020103f
C19001 VDD.t3309 VSS 0.045134f
C19002 VDD.t2033 VSS 0.051441f
C19003 VDD.t1791 VSS 0.020103f
C19004 VDD.t2622 VSS 0.039221f
C19005 VDD.t2416 VSS 0.041192f
C19006 VDD.t2997 VSS 0.049076f
C19007 VDD.t1218 VSS 0.088298f
C19008 VDD.t1787 VSS 0.078178f
C19009 VDD.n2116 VSS 0.121999f
C19010 VDD.n2117 VSS 0.019165f
C19011 VDD.n2118 VSS 0.018088f
C19012 VDD.n2121 VSS 0.016837f
C19013 VDD.n2122 VSS 0.013625f
C19014 VDD.n2127 VSS 0.028241f
C19015 VDD.n2128 VSS 0.013576f
C19016 VDD.n2129 VSS 0.010742f
C19017 VDD.n2130 VSS 0.010413f
C19018 VDD.n2131 VSS 0.011891f
C19019 VDD.n2134 VSS 0.013548f
C19020 VDD.n2135 VSS 0.011852f
C19021 VDD.n2137 VSS 0.013359f
C19022 VDD.n2140 VSS 0.01475f
C19023 VDD.n2144 VSS 0.010788f
C19024 VDD.n2147 VSS 0.014246f
C19025 VDD.n2148 VSS 0.010258f
C19026 VDD.n2149 VSS 0.010392f
C19027 VDD.n2150 VSS 0.118404f
C19028 VDD.n2151 VSS 0.118404f
C19029 VDD.n2157 VSS 0.011115f
C19030 VDD.n2158 VSS 0.015714f
C19031 VDD.n2159 VSS 0.014729f
C19032 VDD.n2160 VSS 0.01408f
C19033 VDD.n2163 VSS 0.011115f
C19034 VDD.n2164 VSS 0.014181f
C19035 VDD.n2165 VSS 0.014295f
C19036 VDD.n2166 VSS 0.015162f
C19037 VDD.n2167 VSS 0.011193f
C19038 VDD.n2168 VSS 0.011509f
C19039 VDD.n2169 VSS 0.014806f
C19040 VDD.n2170 VSS 0.014067f
C19041 VDD.n2171 VSS 0.012133f
C19042 VDD.n2172 VSS 0.010586f
C19043 VDD.n2173 VSS 0.01408f
C19044 VDD.n2174 VSS 0.043882f
C19045 VDD.t3716 VSS 0.061296f
C19046 VDD.t2233 VSS 0.049076f
C19047 VDD.t3558 VSS 0.034097f
C19048 VDD.t1265 VSS 0.039221f
C19049 VDD.t4244 VSS 0.032126f
C19050 VDD.t4242 VSS 0.027002f
C19051 VDD.t2400 VSS 0.022074f
C19052 VDD.t4248 VSS 0.039221f
C19053 VDD.t4246 VSS 0.027002f
C19054 VDD.t4268 VSS 0.022074f
C19055 VDD.t1016 VSS 0.039221f
C19056 VDD.t1012 VSS 0.027002f
C19057 VDD.t1933 VSS 0.022074f
C19058 VDD.t1006 VSS 0.039221f
C19059 VDD.t1004 VSS 0.027002f
C19060 VDD.t2884 VSS 0.022074f
C19061 VDD.t1010 VSS 0.039221f
C19062 VDD.t1018 VSS 0.027002f
C19063 VDD.t4051 VSS 0.022074f
C19064 VDD.t1014 VSS 0.039221f
C19065 VDD.t1008 VSS 0.027002f
C19066 VDD.t1662 VSS 0.038915f
C19067 VDD.n2175 VSS 0.109514f
C19068 VDD.n2187 VSS 0.010992f
C19069 VDD.n2188 VSS 0.010392f
C19070 VDD.n2189 VSS 0.118404f
C19071 VDD.n2190 VSS 0.118404f
C19072 VDD.n2191 VSS 0.010392f
C19073 VDD.n2192 VSS 0.015524f
C19074 VDD.n2193 VSS 0.01408f
C19075 VDD.n2194 VSS 0.01013f
C19076 VDD.n2199 VSS 0.014181f
C19077 VDD.n2200 VSS 0.012648f
C19078 VDD.n2208 VSS 0.010568f
C19079 VDD.n2209 VSS 0.01408f
C19080 VDD.n2210 VSS 0.01013f
C19081 VDD.n2228 VSS 0.012547f
C19082 VDD.n2229 VSS 0.01013f
C19083 VDD.n2246 VSS 0.012547f
C19084 VDD.n2247 VSS 0.01013f
C19085 VDD.n2253 VSS 0.118404f
C19086 VDD.n2254 VSS 0.231769f
C19087 VDD.n2255 VSS 0.010392f
C19088 VDD.n2256 VSS 0.016893f
C19089 VDD.n2257 VSS 0.019165f
C19090 VDD.n2258 VSS 0.01013f
C19091 VDD.n2259 VSS 0.011014f
C19092 VDD.n2261 VSS 0.01408f
C19093 VDD.n2262 VSS 0.015552f
C19094 VDD.n2263 VSS 0.019165f
C19095 VDD.n2264 VSS 0.019165f
C19096 VDD.n2265 VSS 0.019165f
C19097 VDD.n2266 VSS 0.019165f
C19098 VDD.n2267 VSS 0.019165f
C19099 VDD.n2268 VSS 0.019165f
C19100 VDD.n2269 VSS 0.019165f
C19101 VDD.n2270 VSS 0.01013f
C19102 VDD.n2276 VSS 0.011014f
C19103 VDD.n2277 VSS 0.04743f
C19104 VDD.t1401 VSS 0.033112f
C19105 VDD.t2067 VSS 0.044149f
C19106 VDD.t3325 VSS 0.044149f
C19107 VDD.t2378 VSS 0.044149f
C19108 VDD.t2166 VSS 0.044149f
C19109 VDD.t4264 VSS 0.044149f
C19110 VDD.t1863 VSS 0.044149f
C19111 VDD.t3271 VSS 0.044149f
C19112 VDD.t2069 VSS 0.044149f
C19113 VDD.t1521 VSS 0.044149f
C19114 VDD.t1405 VSS 0.044149f
C19115 VDD.t1169 VSS 0.044149f
C19116 VDD.t4253 VSS 0.044149f
C19117 VDD.t2772 VSS 0.044149f
C19118 VDD.t2995 VSS 0.044149f
C19119 VDD.t4003 VSS 0.033112f
C19120 VDD.n2278 VSS 0.036393f
C19121 VDD.n2279 VSS 0.036393f
C19122 VDD.t4055 VSS 0.055186f
C19123 VDD.t3351 VSS 0.055186f
C19124 VDD.t4001 VSS 0.044149f
C19125 VDD.t1341 VSS 0.045528f
C19126 VDD.t2877 VSS 0.036068f
C19127 VDD.t3701 VSS 0.031732f
C19128 VDD.t3386 VSS 0.026213f
C19129 VDD.t3700 VSS 0.044149f
C19130 VDD.t3148 VSS 0.048091f
C19131 VDD.t2017 VSS 0.044149f
C19132 VDD.t2770 VSS 0.044149f
C19133 VDD.t4278 VSS 0.044149f
C19134 VDD.t2205 VSS 0.044149f
C19135 VDD.t3997 VSS 0.044149f
C19136 VDD.t1216 VSS 0.044149f
C19137 VDD.t4255 VSS 0.044149f
C19138 VDD.t2196 VSS 0.033112f
C19139 VDD.n2281 VSS 0.04743f
C19140 VDD.t2585 VSS 0.055186f
C19141 VDD.t1763 VSS 0.044149f
C19142 VDD.t4074 VSS 0.039221f
C19143 VDD.t882 VSS 0.039221f
C19144 VDD.t888 VSS 0.027002f
C19145 VDD.t1205 VSS 0.022074f
C19146 VDD.t886 VSS 0.039221f
C19147 VDD.t884 VSS 0.027002f
C19148 VDD.t3226 VSS 0.022074f
C19149 VDD.t629 VSS 0.039221f
C19150 VDD.t655 VSS 0.027002f
C19151 VDD.t2938 VSS 0.022074f
C19152 VDD.t625 VSS 0.039221f
C19153 VDD.t623 VSS 0.027002f
C19154 VDD.t1851 VSS 0.022074f
C19155 VDD.t653 VSS 0.039221f
C19156 VDD.t665 VSS 0.027002f
C19157 VDD.t4099 VSS 0.022074f
C19158 VDD.t657 VSS 0.039221f
C19159 VDD.t627 VSS 0.027002f
C19160 VDD.t3774 VSS 0.038915f
C19161 VDD.n2287 VSS 0.109514f
C19162 VDD.n2304 VSS 0.01408f
C19163 VDD.n2305 VSS 0.01013f
C19164 VDD.n2313 VSS 0.012648f
C19165 VDD.n2314 VSS 0.010021f
C19166 VDD.n2316 VSS 0.013743f
C19167 VDD.n2318 VSS 0.010568f
C19168 VDD.n2319 VSS 0.01408f
C19169 VDD.n2321 VSS 0.01408f
C19170 VDD.n2322 VSS 0.01013f
C19171 VDD.n2332 VSS 0.231769f
C19172 VDD.n2333 VSS 0.344985f
C19173 VDD.n2334 VSS 0.347695f
C19174 VDD.n2335 VSS 18.7184f
C19175 VDD.n2336 VSS 26.963f
.ends

