* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt cap_mim m4_n120_n120 m4_0_0 VSUBS
X0 m4_0_0 m4_n120_n120 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
C0 m4_0_0 m4_n120_n120 0.414359f
C1 m4_0_0 VSUBS 1.18568f
C2 m4_n120_n120 VSUBS 1.06208f
.ends

.subckt TOP common_bottom top_c2 top_c3 top_c4 top_c5 top_c_dummy top_c1 top_c0
Xcap_mim_0[0|0] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[1|0] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[2|0] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[3|0] common_bottom top_c4 VSUBS cap_mim
Xcap_mim_0[4|0] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[5|0] common_bottom top_c4 VSUBS cap_mim
Xcap_mim_0[6|0] common_bottom top_c4 VSUBS cap_mim
Xcap_mim_0[7|0] common_bottom top_c4 VSUBS cap_mim
Xcap_mim_0[0|1] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[1|1] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[2|1] common_bottom top_c4 VSUBS cap_mim
Xcap_mim_0[3|1] common_bottom m5_n4800_6800 VSUBS cap_mim
Xcap_mim_0[4|1] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[5|1] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[6|1] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[7|1] common_bottom top_c3 VSUBS cap_mim
Xcap_mim_0[0|2] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[1|2] common_bottom top_c3 VSUBS cap_mim
Xcap_mim_0[2|2] common_bottom top_c4 VSUBS cap_mim
Xcap_mim_0[3|2] common_bottom m5_n7400_6800 VSUBS cap_mim
Xcap_mim_0[4|2] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[5|2] common_bottom top_c3 VSUBS cap_mim
Xcap_mim_0[6|2] common_bottom top_c2 VSUBS cap_mim
Xcap_mim_0[7|2] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[0|3] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[1|3] common_bottom top_c4 VSUBS cap_mim
Xcap_mim_0[2|3] common_bottom top_c4 VSUBS cap_mim
Xcap_mim_0[3|3] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[4|3] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[5|3] common_bottom top_c1 VSUBS cap_mim
Xcap_mim_0[6|3] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[7|3] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[0|4] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[1|4] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[2|4] common_bottom top_c1 VSUBS cap_mim
Xcap_mim_0[3|4] common_bottom top_c0 VSUBS cap_mim
Xcap_mim_0[4|4] common_bottom top_c_dummy VSUBS cap_mim
Xcap_mim_0[5|4] common_bottom top_c4 VSUBS cap_mim
Xcap_mim_0[6|4] common_bottom top_c4 VSUBS cap_mim
Xcap_mim_0[7|4] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[0|5] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[1|5] common_bottom top_c2 VSUBS cap_mim
Xcap_mim_0[2|5] common_bottom top_c3 VSUBS cap_mim
Xcap_mim_0[3|5] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[4|5] common_bottom top_c2 VSUBS cap_mim
Xcap_mim_0[5|5] common_bottom top_c4 VSUBS cap_mim
Xcap_mim_0[6|5] common_bottom top_c3 VSUBS cap_mim
Xcap_mim_0[7|5] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[0|6] common_bottom top_c3 VSUBS cap_mim
Xcap_mim_0[1|6] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[2|6] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[3|6] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[4|6] common_bottom top_c3 VSUBS cap_mim
Xcap_mim_0[5|6] common_bottom top_c4 VSUBS cap_mim
Xcap_mim_0[6|6] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[7|6] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[0|7] common_bottom top_c4 VSUBS cap_mim
Xcap_mim_0[1|7] common_bottom top_c4 VSUBS cap_mim
Xcap_mim_0[2|7] common_bottom top_c4 VSUBS cap_mim
Xcap_mim_0[3|7] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[4|7] common_bottom top_c4 VSUBS cap_mim
Xcap_mim_0[5|7] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[6|7] common_bottom top_c5 VSUBS cap_mim
Xcap_mim_0[7|7] common_bottom top_c5 VSUBS cap_mim
C0 top_c1 top_c_dummy 0.013909f
C1 top_c0 top_c1 2.053814f
C2 top_c4 common_bottom 20.381252f
C3 top_c_dummy top_c2 2.017989f
C4 top_c3 top_c4 2.710395f
C5 top_c0 top_c2 0.02726f
C6 top_c5 common_bottom 41.545517f
C7 top_c1 top_c2 0.051003f
C8 top_c3 top_c5 2.307618f
C9 m5_n7400_6800 top_c2 0.200803f
C10 top_c4 top_c5 5.341128f
C11 top_c_dummy common_bottom 1.713993f
C12 top_c0 common_bottom 1.428327f
C13 top_c3 top_c_dummy 0.004478f
C14 top_c3 top_c0 5.04e-19
C15 top_c1 common_bottom 2.684169f
C16 m5_n7400_6800 m5_n4800_6800 0.22972f
C17 top_c3 top_c1 5.04e-19
C18 top_c2 common_bottom 6.281751f
C19 top_c4 top_c_dummy 0.362575f
C20 m5_n7400_6800 common_bottom 0.497373f
C21 top_c4 top_c0 0.208334f
C22 top_c3 top_c2 1.055012f
C23 top_c3 m5_n7400_6800 0.038421f
C24 top_c4 top_c1 0.381888f
C25 top_c5 top_c_dummy 0.295218f
C26 top_c5 top_c0 0.439582f
C27 m5_n4800_6800 common_bottom 0.532008f
C28 top_c4 top_c2 0.285824f
C29 top_c5 top_c1 0.622374f
C30 top_c3 m5_n4800_6800 0.235662f
C31 top_c5 top_c2 1.279418f
C32 top_c5 m5_n7400_6800 0.11486f
C33 top_c3 common_bottom 8.641127f
C34 top_c0 top_c_dummy 0.089269f
C35 top_c4 m5_n4800_6800 0.056913f
C36 top_c5 VSUBS 62.147964f
C37 top_c4 VSUBS 38.041428f
C38 common_bottom VSUBS 0.118965p
C39 top_c_dummy VSUBS 3.679576f
C40 top_c0 VSUBS 4.36327f
C41 top_c1 VSUBS 6.20843f
C42 top_c2 VSUBS 12.04523f
C43 m5_n7400_6800 VSUBS 1.14708f
C44 top_c3 VSUBS 22.510658f
C45 m5_n4800_6800 VSUBS 1.305221f
.ends

