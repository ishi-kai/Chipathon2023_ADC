* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt TOP top_c4 top_c3 top_c2 top_c_dummy top_c0 top_c1 common_bottom top_c5
X0 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X1 top_c3 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X2 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X3 top_c3 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X4 top_c4 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X5 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X6 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X7 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X8 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X9 top_c0 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X10 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X11 top_c3 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X12 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X13 top_c3 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X14 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X15 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X16 top_c2 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X17 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X18 top_c4 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X19 top_c3 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X20 top_c4 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X21 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X22 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X23 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X24 top_c4 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X25 top_c4 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X26 top_c4 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X27 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X28 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X29 top_c4 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X30 top_c4 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X31 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X32 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X33 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X34 top_c4 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X35 top_c2 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X36 top_c4 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X37 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X38 top_c_dummy common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X39 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X40 top_c2 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X41 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X42 top_c1 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X43 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X44 top_c4 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X45 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X46 top_c1 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X47 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X48 top_c4 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X49 top_c4 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X50 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X51 top_c3 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X52 top_c4 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X53 top_c4 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X54 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X55 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X56 top_c3 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X57 top_c4 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X58 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X59 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X60 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X61 top_c3 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X62 top_c2 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X63 top_c5 common_bottom cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
C0 m3_13080_37400 top_c4 0.17689f
C1 top_c0 top_c4 0.344447f
C2 m3_n1920_37400 top_c4 3.57873f
C3 m3_13080_37400 top_c3 3.68826f
C4 m3_n1920_37400 top_c3 0.283216f
C5 top_c2 top_c_dummy 3.90557f
C6 top_c0 top_c3 0.07203f
C7 m3_9600_37600 common_bottom 1.11158f
C8 m3_9600_37600 top_c4 0.334345f
C9 m3_9600_37600 top_c3 0.031939f
C10 top_c2 top_c5 2.51643f
C11 m3_1080_37400 top_c5 0.499167f
C12 common_bottom m3_16080_37400 1.11115f
C13 top_c4 m3_16080_37400 4.00191f
C14 m3_16080_37400 top_c3 0.023466f
C15 top_c1 top_c2 0.113754f
C16 top_c_dummy common_bottom 2.16056f
C17 top_c_dummy top_c4 0.557255f
C18 top_c_dummy top_c3 0.103688f
C19 top_c2 m3_1080_37400 0.31178f
C20 common_bottom top_c5 34.3926f
C21 top_c4 top_c5 10.3785f
C22 top_c3 top_c5 3.25187f
C23 top_c1 common_bottom 3.26961f
C24 top_c1 top_c4 0.488545f
C25 top_c1 top_c3 0.35918f
C26 top_c2 common_bottom 6.95875f
C27 m3_1080_37400 common_bottom 1.11094f
C28 top_c2 top_c4 0.834243f
C29 m3_1080_37400 top_c4 0.175599f
C30 top_c_dummy top_c0 0.470294f
C31 top_c2 top_c3 3.36078f
C32 m3_1080_37400 top_c3 3.70845f
C33 m3_13080_37400 top_c5 0.804673f
C34 m3_n1920_37400 top_c5 0.833773f
C35 top_c0 top_c5 0.872246f
C36 m3_9600_37600 top_c5 0.782903f
C37 top_c1 top_c0 3.94932f
C38 top_c1 m3_9600_37600 0.15589f
C39 common_bottom top_c4 17.7895f
C40 common_bottom top_c3 10.7252f
C41 top_c4 top_c3 5.28718f
C42 m3_16080_37400 top_c5 0.68244f
C43 top_c2 m3_13080_37400 0.0295f
C44 top_c2 top_c0 0.097925f
C45 top_c2 m3_9600_37600 3.35976f
C46 top_c_dummy top_c5 0.696513f
C47 top_c1 top_c_dummy 0.171719f
C48 common_bottom m3_13080_37400 1.11094f
C49 m3_n1920_37400 common_bottom 1.11032f
C50 top_c1 top_c5 1.32165f
C51 top_c0 common_bottom 2.17708f
C52 common_bottom VSUBS 80.762f
C53 top_c1 VSUBS 9.66846f
C54 top_c0 VSUBS 7.34352f
C55 top_c_dummy VSUBS 7.33815f
C56 top_c2 VSUBS 19.648699f
C57 top_c3 VSUBS 28.811598f
C58 top_c4 VSUBS 45.077602f
C59 top_c5 VSUBS 85.211205f
C60 m3_16080_37400 VSUBS 4.82137f $ **FLOATING
C61 m3_13080_37400 VSUBS 4.82148f $ **FLOATING
C62 m3_9600_37600 VSUBS 4.77941f $ **FLOATING
C63 m3_1080_37400 VSUBS 4.82141f $ **FLOATING
C64 m3_n1920_37400 VSUBS 4.82137f $ **FLOATING
.ends

