* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt TOP S R VDD GND Qn Q
X0 Q.t0 Qn.t3 GND.t7 GND.t6 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X1 VDD.t1 R.t0 a_2894_1087 VDD.t0 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X2 GND.t5 a_85_1225 Qn.t1 GND.t4 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X3 Q.t2 a_2894_1087 GND.t9 GND.t8 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X4 GND.t11 R.t1 a_2894_1087 GND.t10 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X5 a_85_1225 S.t0 VDD.t7 VDD.t6 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X6 VDD.t3 Q.t3 Qn.t2 VDD.t2 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X7 a_85_1225 S.t1 GND.t3 GND.t2 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X8 GND.t1 Q.t4 Qn.t0 GND.t0 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X9 Q.t1 Qn.t4 VDD.t5 VDD.t4 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
R0 Qn Qn.t4 56.0856
R1 Qn.n1 Qn.t3 55.9719
R2 Qn.n2 Qn.t1 4.35469
R3 Qn.n1 Qn.n0 3.18045
R4 Qn.n0 Qn.t2 3.0207
R5 Qn.n0 Qn.t0 2.1605
R6 Qn.n2 Qn.n1 0.068
R7 Qn Qn.n2 0.0573421
R8 GND.n12 GND.n3 31486
R9 GND.n13 GND.n12 30891.4
R10 GND.n12 GND.n11 9378.27
R11 GND.t4 GND.t2 1731.97
R12 GND.t10 GND.t8 1592.53
R13 GND.n11 GND.t0 1534.44
R14 GND.n11 GND.t6 1534.44
R15 GND.n5 GND.t10 856.457
R16 GND.t0 GND.n10 854.365
R17 GND.t6 GND.n2 854.365
R18 GND.n17 GND.t2 851.1
R19 GND.n14 GND.n2 795.389
R20 GND.n10 GND.n4 792.851
R21 GND.n14 GND.n13 719.958
R22 GND.n4 GND.n3 649.317
R23 GND.t8 GND.n3 205.048
R24 GND.n13 GND.t4 129.049
R25 GND.n17 GND.n16 5.86657
R26 GND.n7 GND.n5 5.78782
R27 GND.n7 GND.n6 4.5005
R28 GND.n9 GND.n8 4.5005
R29 GND.n1 GND.n0 4.5005
R30 GND.n16 GND.n15 4.5005
R31 GND.n6 GND.t9 2.17407
R32 GND.n9 GND.t1 2.17389
R33 GND.n5 GND.t11 2.17352
R34 GND.n1 GND.t7 2.17333
R35 GND.n15 GND.t5 2.17314
R36 GND GND.t3 2.16794
R37 GND.n15 GND.n14 2.09426
R38 GND.n2 GND.n1 2.09407
R39 GND.n10 GND.n9 2.09352
R40 GND.n6 GND.n4 2.09333
R41 GND.n8 GND.n0 1.97889
R42 GND.n16 GND.n0 0.572643
R43 GND.n8 GND.n7 0.558179
R44 GND GND.n17 0.00793802
R45 Q.n2 Q.t4 56.0619
R46 Q.n1 Q.t3 55.9719
R47 Q.n2 Q.t2 4.38208
R48 Q.n1 Q.n0 3.62303
R49 Q.n0 Q.t0 3.0907
R50 Q.n0 Q.t1 2.0905
R51 Q Q.n1 0.108263
R52 Q Q.n2 0.0407632
R53 R R.t0 56.1318
R54 R R.t1 56.0501
R55 VDD.n0 VDD.t0 311.147
R56 VDD.n1 VDD.t2 311.146
R57 VDD.n5 VDD.t6 311.132
R58 VDD.n3 VDD.t4 311.132
R59 VDD.n5 VDD.n4 6.45318
R60 VDD.n2 VDD.n0 6.38568
R61 VDD.n4 VDD.n3 4.50293
R62 VDD.n2 VDD.n1 4.5005
R63 VDD.n1 VDD.t3 2.10463
R64 VDD.n0 VDD.t1 2.10445
R65 VDD.n5 VDD.t7 2.0905
R66 VDD.n3 VDD.t5 2.0905
R67 VDD.n4 VDD.n2 2.01104
R68 VDD VDD.n5 0.0540135
R69 S S.t0 56.0986
R70 S S.t1 56.0832
C0 Qn a_85_1225 0.291767f
C1 Qn Q 1.62575f
C2 R a_2894_1087 0.16834f
C3 Q a_2894_1087 0.378711f
C4 Qn VDD 0.403238f
C5 VDD a_85_1225 0.347733f
C6 a_2894_1087 VDD 0.349789f
C7 S a_85_1225 0.167843f
C8 R VDD 0.174505f
C9 Q VDD 1.17919f
C10 S VDD 0.174547f
C11 R GND 0.347354f
C12 Q GND 1.54705f
C13 Qn GND 2.3216f
C14 S GND 0.348389f
C15 VDD GND 8.457769f
C16 a_2894_1087 GND 0.83604f
C17 a_85_1225 GND 0.875087f
.ends

