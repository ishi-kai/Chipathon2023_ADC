* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt TOP top_c5 top_c3 top_c2 top_c4 top_c0 top_c1 top_c_dummy common_bottom
X0 top_c5.t0 common_bottom.t56 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X1 top_c3.t0 common_bottom.t13 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X2 top_c5.t1 common_bottom.t55 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X3 top_c3.t1 common_bottom.t61 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X4 top_c4.t0 common_bottom.t21 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X5 top_c5.t2 common_bottom.t54 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X6 top_c5.t3 common_bottom.t53 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X7 top_c5.t4 common_bottom.t52 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X8 top_c5.t5 common_bottom.t51 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X9 top_c0.t0 common_bottom.t14 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X10 top_c5.t6 common_bottom.t50 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X11 top_c3.t2 common_bottom.t2 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X12 top_c5.t7 common_bottom.t49 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X13 top_c3.t3 common_bottom.t1 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X14 top_c5.t8 common_bottom.t48 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X15 top_c5.t9 common_bottom.t47 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X16 top_c2.t0 common_bottom.t11 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X17 top_c5.t10 common_bottom.t46 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X18 top_c4.t1 common_bottom.t9 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X19 top_c3.t4 common_bottom.t7 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X20 top_c4.t2 common_bottom.t16 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X21 top_c5.t11 common_bottom.t45 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X22 top_c5.t12 common_bottom.t44 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X23 top_c5.t13 common_bottom.t43 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X24 top_c4.t3 common_bottom.t62 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X25 top_c4.t4 common_bottom.t15 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X26 top_c4.t5 common_bottom.t59 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X27 top_c5.t14 common_bottom.t42 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X28 top_c5.t15 common_bottom.t41 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X29 top_c4.t6 common_bottom.t23 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X30 top_c4.t7 common_bottom.t63 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X31 top_c5.t16 common_bottom.t40 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X32 top_c5.t17 common_bottom.t39 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X33 top_c5.t18 common_bottom.t38 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X34 top_c4.t8 common_bottom.t5 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X35 top_c2.t1 common_bottom.t0 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X36 top_c4.t9 common_bottom.t20 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X37 top_c5.t19 common_bottom.t37 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X38 top_c_dummy.t0 common_bottom.t12 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X39 top_c5.t20 common_bottom.t36 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X40 top_c2.t2 common_bottom.t60 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X41 top_c5.t21 common_bottom.t35 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X42 top_c0.t1 common_bottom.t3 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X43 top_c5.t22 common_bottom.t34 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X44 top_c4.t10 common_bottom.t58 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X45 top_c5.t23 common_bottom.t33 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X46 top_c1.t0 common_bottom.t19 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X47 top_c5.t24 common_bottom.t32 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X48 top_c4.t11 common_bottom.t22 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X49 top_c4.t12 common_bottom.t57 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X50 top_c5.t25 common_bottom.t31 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X51 top_c3.t5 common_bottom.t17 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X52 top_c4.t13 common_bottom.t6 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X53 top_c4.t14 common_bottom.t8 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X54 top_c5.t26 common_bottom.t30 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X55 top_c5.t27 common_bottom.t29 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X56 top_c3.t6 common_bottom.t10 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X57 top_c4.t15 common_bottom.t4 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X58 top_c5.t28 common_bottom.t28 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X59 top_c5.t29 common_bottom.t27 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X60 top_c5.t30 common_bottom.t26 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X61 top_c3.t7 common_bottom.t24 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X62 top_c2.t3 common_bottom.t18 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X63 top_c5.t31 common_bottom.t25 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
R0 top_c5.n198 top_c5.n197 39.854
R1 top_c5.n183 top_c5.n182 5.2655
R2 top_c5.n56 top_c5.n55 5.2655
R3 top_c5.n192 top_c5.n183 4.5675
R4 top_c5.n188 top_c5.n112 4.5675
R5 top_c5.n59 top_c5.n56 4.5675
R6 top_c5.n62 top_c5.n61 4.5675
R7 top_c5.n195 top_c5.n100 4.5005
R8 top_c5.n196 top_c5.n195 4.5005
R9 top_c5.n159 top_c5.n119 4.5005
R10 top_c5.n155 top_c5.n119 4.5005
R11 top_c5.n145 top_c5.n126 4.5005
R12 top_c5.n141 top_c5.n126 4.5005
R13 top_c5.n138 top_c5.n117 4.5005
R14 top_c5.n134 top_c5.n117 4.5005
R15 top_c5.n180 top_c5.n115 4.5005
R16 top_c5.n181 top_c5.n180 4.5005
R17 top_c5.n152 top_c5.n123 4.5005
R18 top_c5.n148 top_c5.n123 4.5005
R19 top_c5.n160 top_c5.n159 4.5005
R20 top_c5.n158 top_c5.n120 4.5005
R21 top_c5.n156 top_c5.n121 4.5005
R22 top_c5.n155 top_c5.n154 4.5005
R23 top_c5.n153 top_c5.n152 4.5005
R24 top_c5.n151 top_c5.n122 4.5005
R25 top_c5.n149 top_c5.n124 4.5005
R26 top_c5.n148 top_c5.n147 4.5005
R27 top_c5.n146 top_c5.n145 4.5005
R28 top_c5.n144 top_c5.n125 4.5005
R29 top_c5.n142 top_c5.n127 4.5005
R30 top_c5.n141 top_c5.n140 4.5005
R31 top_c5.n139 top_c5.n138 4.5005
R32 top_c5.n137 top_c5.n128 4.5005
R33 top_c5.n135 top_c5.n129 4.5005
R34 top_c5.n134 top_c5.n133 4.5005
R35 top_c5.n132 top_c5.n115 4.5005
R36 top_c5.n131 top_c5.n130 4.5005
R37 top_c5.n114 top_c5.n113 4.5005
R38 top_c5.n182 top_c5.n181 4.5005
R39 top_c5.n191 top_c5.n190 4.5005
R40 top_c5.n189 top_c5.n184 4.5005
R41 top_c5.n187 top_c5.n100 4.5005
R42 top_c5.n186 top_c5.n185 4.5005
R43 top_c5.n99 top_c5.n98 4.5005
R44 top_c5.n197 top_c5.n196 4.5005
R45 top_c5.n67 top_c5.n34 4.5005
R46 top_c5.n68 top_c5.n67 4.5005
R47 top_c5.n81 top_c5.n10 4.5005
R48 top_c5.n82 top_c5.n81 4.5005
R49 top_c5.n74 top_c5.n13 4.5005
R50 top_c5.n75 top_c5.n74 4.5005
R51 top_c5.n95 top_c5.n3 4.5005
R52 top_c5.n96 top_c5.n95 4.5005
R53 top_c5.n88 top_c5.n6 4.5005
R54 top_c5.n89 top_c5.n88 4.5005
R55 top_c5.n53 top_c5.n48 4.5005
R56 top_c5.n54 top_c5.n53 4.5005
R57 top_c5.n49 top_c5.n48 4.5005
R58 top_c5.n51 top_c5.n50 4.5005
R59 top_c5.n38 top_c5.n37 4.5005
R60 top_c5.n55 top_c5.n54 4.5005
R61 top_c5.n58 top_c5.n57 4.5005
R62 top_c5.n36 top_c5.n35 4.5005
R63 top_c5.n63 top_c5.n34 4.5005
R64 top_c5.n65 top_c5.n64 4.5005
R65 top_c5.n15 top_c5.n14 4.5005
R66 top_c5.n69 top_c5.n68 4.5005
R67 top_c5.n70 top_c5.n13 4.5005
R68 top_c5.n72 top_c5.n71 4.5005
R69 top_c5.n12 top_c5.n11 4.5005
R70 top_c5.n76 top_c5.n75 4.5005
R71 top_c5.n77 top_c5.n10 4.5005
R72 top_c5.n79 top_c5.n78 4.5005
R73 top_c5.n8 top_c5.n7 4.5005
R74 top_c5.n83 top_c5.n82 4.5005
R75 top_c5.n84 top_c5.n6 4.5005
R76 top_c5.n86 top_c5.n85 4.5005
R77 top_c5.n5 top_c5.n4 4.5005
R78 top_c5.n90 top_c5.n89 4.5005
R79 top_c5.n91 top_c5.n3 4.5005
R80 top_c5.n93 top_c5.n92 4.5005
R81 top_c5.n1 top_c5.n0 4.5005
R82 top_c5.n97 top_c5.n96 4.5005
R83 top_c5.n49 top_c5.n47 3.09683
R84 top_c5.n161 top_c5.n160 3.09583
R85 top_c5.n195 top_c5.n101 2.21775
R86 top_c5.n193 top_c5.n192 2.21775
R87 top_c5.n193 top_c5.n112 2.21775
R88 top_c5.n157 top_c5.n119 2.21775
R89 top_c5.n143 top_c5.n126 2.21775
R90 top_c5.n136 top_c5.n117 2.21775
R91 top_c5.n180 top_c5.n116 2.21775
R92 top_c5.n150 top_c5.n123 2.21775
R93 top_c5.n67 top_c5.n66 2.21775
R94 top_c5.n81 top_c5.n80 2.21775
R95 top_c5.n74 top_c5.n73 2.21775
R96 top_c5.n95 top_c5.n94 2.21775
R97 top_c5.n88 top_c5.n87 2.21775
R98 top_c5.n60 top_c5.n59 2.21775
R99 top_c5.n61 top_c5.n60 2.21775
R100 top_c5.n53 top_c5.n52 2.21775
R101 top_c5.n140 top_c5.n139 1.8905
R102 top_c5.n84 top_c5.n83 1.8905
R103 top_c5.n154 top_c5.n153 1.88938
R104 top_c5.n70 top_c5.n69 1.88938
R105 top_c5.n198 top_c5.n97 1.6893
R106 top_c5.n105 top_c5.n103 0.988357
R107 top_c5.n103 top_c5.n102 0.988357
R108 top_c5.n166 top_c5.n165 0.988357
R109 top_c5.n168 top_c5.n165 0.988357
R110 top_c5.n171 top_c5.n164 0.988357
R111 top_c5.n20 top_c5.n19 0.988357
R112 top_c5.n22 top_c5.n19 0.988357
R113 top_c5.n25 top_c5.n18 0.988357
R114 top_c5.n27 top_c5.n18 0.988357
R115 top_c5.n30 top_c5.n16 0.988357
R116 top_c5.n40 top_c5.n39 0.988357
R117 top_c5.n42 top_c5.n40 0.988357
R118 top_c5.n173 top_c5.n164 0.988261
R119 top_c5.n177 top_c5.n176 0.987576
R120 top_c5.n176 top_c5.n174 0.960525
R121 top_c5.n110 top_c5.n102 0.9605
R122 top_c5.n108 top_c5.n105 0.9605
R123 top_c5.n178 top_c5.n118 0.9605
R124 top_c5.n162 top_c5.n118 0.9605
R125 top_c5.n32 top_c5.n17 0.9605
R126 top_c5.n30 top_c5.n29 0.9605
R127 top_c5.n43 top_c5.n42 0.9605
R128 top_c5.n45 top_c5.n39 0.9605
R129 top_c5.n33 top_c5.n32 0.9599
R130 top_c5.n147 top_c5.n146 0.676625
R131 top_c5.n63 top_c5.n62 0.676625
R132 top_c5.n133 top_c5.n132 0.6755
R133 top_c5.n188 top_c5.n187 0.6755
R134 top_c5.n77 top_c5.n76 0.6755
R135 top_c5.n91 top_c5.n90 0.6755
R136 top_c5.n166 top_c5.t2 0.60448
R137 top_c5.n20 top_c5.t5 0.60448
R138 top_c5.n43 top_c5.t18 0.60448
R139 top_c5.n106 top_c5.t25 0.586765
R140 top_c5.n170 top_c5.n169 0.5405
R141 top_c5.n24 top_c5.n23 0.5405
R142 top_c5.n107 top_c5.n106 0.526689
R143 top_c5.n108 top_c5.n107 0.512643
R144 top_c5.n171 top_c5.n170 0.512643
R145 top_c5.n25 top_c5.n24 0.512643
R146 top_c5.n111 top_c5.n110 0.512643
R147 top_c5.n169 top_c5.n168 0.512643
R148 top_c5.n23 top_c5.n22 0.512643
R149 top_c5.n46 top_c5.n45 0.512643
R150 top_c5 top_c5.n198 0.494559
R151 top_c5.n174 top_c5.n173 0.484786
R152 top_c5.n29 top_c5.n27 0.484786
R153 top_c5.n185 top_c5.n100 0.1355
R154 top_c5.n196 top_c5.n99 0.1355
R155 top_c5.n191 top_c5.n184 0.1355
R156 top_c5.n159 top_c5.n158 0.1355
R157 top_c5.n156 top_c5.n155 0.1355
R158 top_c5.n145 top_c5.n144 0.1355
R159 top_c5.n142 top_c5.n141 0.1355
R160 top_c5.n130 top_c5.n115 0.1355
R161 top_c5.n181 top_c5.n114 0.1355
R162 top_c5.n138 top_c5.n137 0.1355
R163 top_c5.n135 top_c5.n134 0.1355
R164 top_c5.n152 top_c5.n151 0.1355
R165 top_c5.n149 top_c5.n148 0.1355
R166 top_c5.n160 top_c5.n120 0.1355
R167 top_c5.n121 top_c5.n120 0.1355
R168 top_c5.n154 top_c5.n121 0.1355
R169 top_c5.n153 top_c5.n122 0.1355
R170 top_c5.n124 top_c5.n122 0.1355
R171 top_c5.n147 top_c5.n124 0.1355
R172 top_c5.n146 top_c5.n125 0.1355
R173 top_c5.n127 top_c5.n125 0.1355
R174 top_c5.n140 top_c5.n127 0.1355
R175 top_c5.n139 top_c5.n128 0.1355
R176 top_c5.n129 top_c5.n128 0.1355
R177 top_c5.n133 top_c5.n129 0.1355
R178 top_c5.n132 top_c5.n131 0.1355
R179 top_c5.n131 top_c5.n113 0.1355
R180 top_c5.n182 top_c5.n113 0.1355
R181 top_c5.n190 top_c5.n183 0.1355
R182 top_c5.n190 top_c5.n189 0.1355
R183 top_c5.n189 top_c5.n188 0.1355
R184 top_c5.n187 top_c5.n186 0.1355
R185 top_c5.n186 top_c5.n98 0.1355
R186 top_c5.n197 top_c5.n98 0.1355
R187 top_c5.n65 top_c5.n34 0.1355
R188 top_c5.n68 top_c5.n15 0.1355
R189 top_c5.n72 top_c5.n13 0.1355
R190 top_c5.n75 top_c5.n12 0.1355
R191 top_c5.n79 top_c5.n10 0.1355
R192 top_c5.n82 top_c5.n8 0.1355
R193 top_c5.n86 top_c5.n6 0.1355
R194 top_c5.n89 top_c5.n5 0.1355
R195 top_c5.n93 top_c5.n3 0.1355
R196 top_c5.n96 top_c5.n1 0.1355
R197 top_c5.n58 top_c5.n36 0.1355
R198 top_c5.n51 top_c5.n48 0.1355
R199 top_c5.n54 top_c5.n38 0.1355
R200 top_c5.n50 top_c5.n49 0.1355
R201 top_c5.n50 top_c5.n37 0.1355
R202 top_c5.n55 top_c5.n37 0.1355
R203 top_c5.n57 top_c5.n56 0.1355
R204 top_c5.n57 top_c5.n35 0.1355
R205 top_c5.n62 top_c5.n35 0.1355
R206 top_c5.n64 top_c5.n63 0.1355
R207 top_c5.n64 top_c5.n14 0.1355
R208 top_c5.n69 top_c5.n14 0.1355
R209 top_c5.n71 top_c5.n70 0.1355
R210 top_c5.n71 top_c5.n11 0.1355
R211 top_c5.n76 top_c5.n11 0.1355
R212 top_c5.n78 top_c5.n77 0.1355
R213 top_c5.n78 top_c5.n7 0.1355
R214 top_c5.n83 top_c5.n7 0.1355
R215 top_c5.n85 top_c5.n84 0.1355
R216 top_c5.n85 top_c5.n4 0.1355
R217 top_c5.n90 top_c5.n4 0.1355
R218 top_c5.n92 top_c5.n91 0.1355
R219 top_c5.n92 top_c5.n0 0.1355
R220 top_c5.n97 top_c5.n0 0.1355
R221 top_c5.n106 top_c5.t10 0.106765
R222 top_c5.n107 top_c5.t23 0.0923367
R223 top_c5.n103 top_c5.t11 0.0923367
R224 top_c5.n104 top_c5.t26 0.0923367
R225 top_c5.n109 top_c5.t12 0.0923367
R226 top_c5.n111 top_c5.t29 0.0923367
R227 top_c5.n165 top_c5.t8 0.0923367
R228 top_c5.n167 top_c5.t24 0.0923367
R229 top_c5.n169 top_c5.t13 0.0923367
R230 top_c5.n170 top_c5.t27 0.0923367
R231 top_c5.n164 top_c5.t28 0.0923367
R232 top_c5.n172 top_c5.t14 0.0923367
R233 top_c5.n177 top_c5.t30 0.0923367
R234 top_c5.n175 top_c5.t16 0.0923367
R235 top_c5.n163 top_c5.t0 0.0923367
R236 top_c5.n19 top_c5.t7 0.0923367
R237 top_c5.n21 top_c5.t22 0.0923367
R238 top_c5.n23 top_c5.t1 0.0923367
R239 top_c5.n24 top_c5.t15 0.0923367
R240 top_c5.n18 top_c5.t31 0.0923367
R241 top_c5.n26 top_c5.t17 0.0923367
R242 top_c5.n28 top_c5.t4 0.0923367
R243 top_c5.n31 top_c5.t20 0.0923367
R244 top_c5.n16 top_c5.t6 0.0923367
R245 top_c5.n40 top_c5.t21 0.0923367
R246 top_c5.n41 top_c5.t3 0.0923367
R247 top_c5.n44 top_c5.t19 0.0923367
R248 top_c5.n46 top_c5.t9 0.0923367
R249 top_c5.n101 top_c5.n99 0.0675025
R250 top_c5.n185 top_c5.n101 0.0675025
R251 top_c5.n184 top_c5.n112 0.0675025
R252 top_c5.n192 top_c5.n191 0.0675025
R253 top_c5.n157 top_c5.n156 0.0675025
R254 top_c5.n158 top_c5.n157 0.0675025
R255 top_c5.n143 top_c5.n142 0.0675025
R256 top_c5.n144 top_c5.n143 0.0675025
R257 top_c5.n116 top_c5.n114 0.0675025
R258 top_c5.n136 top_c5.n135 0.0675025
R259 top_c5.n137 top_c5.n136 0.0675025
R260 top_c5.n130 top_c5.n116 0.0675025
R261 top_c5.n150 top_c5.n149 0.0675025
R262 top_c5.n151 top_c5.n150 0.0675025
R263 top_c5.n66 top_c5.n15 0.0675025
R264 top_c5.n66 top_c5.n65 0.0675025
R265 top_c5.n73 top_c5.n12 0.0675025
R266 top_c5.n80 top_c5.n8 0.0675025
R267 top_c5.n80 top_c5.n79 0.0675025
R268 top_c5.n73 top_c5.n72 0.0675025
R269 top_c5.n87 top_c5.n5 0.0675025
R270 top_c5.n94 top_c5.n1 0.0675025
R271 top_c5.n94 top_c5.n93 0.0675025
R272 top_c5.n87 top_c5.n86 0.0675025
R273 top_c5.n61 top_c5.n36 0.0675025
R274 top_c5.n59 top_c5.n58 0.0675025
R275 top_c5.n52 top_c5.n38 0.0675025
R276 top_c5.n52 top_c5.n51 0.0675025
R277 top_c5.n195 top_c5.n194 0.0557273
R278 top_c5.n194 top_c5.n193 0.0557273
R279 top_c5.n161 top_c5.n119 0.0557273
R280 top_c5.n126 top_c5.n118 0.0557273
R281 top_c5.n179 top_c5.n117 0.0557273
R282 top_c5.n180 top_c5.n179 0.0557273
R283 top_c5.n123 top_c5.n118 0.0557273
R284 top_c5.n67 top_c5.n33 0.0557273
R285 top_c5.n81 top_c5.n9 0.0557273
R286 top_c5.n74 top_c5.n9 0.0557273
R287 top_c5.n95 top_c5.n2 0.0557273
R288 top_c5.n88 top_c5.n2 0.0557273
R289 top_c5.n60 top_c5.n33 0.0557273
R290 top_c5.n53 top_c5.n47 0.0557273
R291 top_c5.n194 top_c5.n111 0.0305
R292 top_c5.n47 top_c5.n46 0.0305
R293 top_c5.n176 top_c5.n175 0.029221
R294 top_c5.n33 top_c5.n16 0.0288259
R295 top_c5.n104 top_c5.n102 0.0283571
R296 top_c5.n105 top_c5.n104 0.0283571
R297 top_c5.n110 top_c5.n109 0.0283571
R298 top_c5.n109 top_c5.n108 0.0283571
R299 top_c5.n168 top_c5.n167 0.0283571
R300 top_c5.n167 top_c5.n166 0.0283571
R301 top_c5.n173 top_c5.n172 0.0283571
R302 top_c5.n172 top_c5.n171 0.0283571
R303 top_c5.n178 top_c5.n177 0.0283571
R304 top_c5.n175 top_c5.n118 0.0283571
R305 top_c5.n163 top_c5.n162 0.0283571
R306 top_c5.n174 top_c5.n163 0.0283571
R307 top_c5.n21 top_c5.n20 0.0283571
R308 top_c5.n22 top_c5.n21 0.0283571
R309 top_c5.n26 top_c5.n25 0.0283571
R310 top_c5.n27 top_c5.n26 0.0283571
R311 top_c5.n29 top_c5.n28 0.0283571
R312 top_c5.n28 top_c5.n17 0.0283571
R313 top_c5.n31 top_c5.n30 0.0283571
R314 top_c5.n32 top_c5.n31 0.0283571
R315 top_c5.n42 top_c5.n41 0.0283571
R316 top_c5.n41 top_c5.n39 0.0283571
R317 top_c5.n44 top_c5.n43 0.0283571
R318 top_c5.n45 top_c5.n44 0.0283571
R319 top_c5.n179 top_c5.n178 0.00264286
R320 top_c5.n162 top_c5.n161 0.00264286
R321 top_c5.n17 top_c5.n2 0.00264286
R322 top_c5.n32 top_c5.n9 0.00264286
R323 common_bottom common_bottom.t15 3.05781
R324 common_bottom.t6 common_bottom.t1 1.23983
R325 common_bottom.t1 common_bottom.t54 1.23983
R326 common_bottom.t54 common_bottom.t32 1.23983
R327 common_bottom.t32 common_bottom.t43 1.23983
R328 common_bottom.t29 common_bottom.t43 1.23983
R329 common_bottom.t42 common_bottom.t29 1.23983
R330 common_bottom.t17 common_bottom.t51 1.23216
R331 common_bottom.t60 common_bottom.t45 1.23216
R332 common_bottom.t30 common_bottom.t2 1.23216
R333 common_bottom.t44 common_bottom.t33 1.23216
R334 common_bottom.t10 common_bottom.t11 1.23216
R335 common_bottom.t62 common_bottom.t57 1.23216
R336 common_bottom.t7 common_bottom.t28 1.23216
R337 common_bottom.t51 common_bottom.t34 1.23216
R338 common_bottom.t34 common_bottom.t55 1.23216
R339 common_bottom.t49 common_bottom.t20 1.23216
R340 common_bottom.t19 common_bottom.t21 1.23216
R341 common_bottom.t46 common_bottom.t12 1.23216
R342 common_bottom.t31 common_bottom.t14 1.23216
R343 common_bottom.t8 common_bottom.t48 1.23216
R344 common_bottom.t48 common_bottom.t0 1.23216
R345 common_bottom.t41 common_bottom.t39 1.23216
R346 common_bottom.t39 common_bottom.t52 1.23216
R347 common_bottom.t36 common_bottom.t25 1.23216
R348 common_bottom.t50 common_bottom.t5 1.23216
R349 common_bottom.t58 common_bottom.t61 1.23216
R350 common_bottom.t47 common_bottom.t37 1.23216
R351 common_bottom.t22 common_bottom.t53 1.23216
R352 common_bottom.t9 common_bottom.t35 1.23216
R353 common_bottom.t56 common_bottom.t42 1.23216
R354 common_bottom.t17 common_bottom.t45 1.2245
R355 common_bottom.t30 common_bottom.t45 1.2245
R356 common_bottom.t30 common_bottom.t44 1.2245
R357 common_bottom.t44 common_bottom.t10 1.2245
R358 common_bottom.t10 common_bottom.t62 1.2245
R359 common_bottom.t28 common_bottom.t62 1.2245
R360 common_bottom.t28 common_bottom.t42 1.2245
R361 common_bottom.t20 common_bottom.t55 1.2245
R362 common_bottom.t21 common_bottom.t20 1.2245
R363 common_bottom.t12 common_bottom.t21 1.2245
R364 common_bottom.t14 common_bottom.t12 1.2245
R365 common_bottom.t3 common_bottom.t14 1.2245
R366 common_bottom.t7 common_bottom.t29 1.2245
R367 common_bottom.t7 common_bottom.t57 1.2245
R368 common_bottom.t57 common_bottom.t11 1.2245
R369 common_bottom.t11 common_bottom.t33 1.2245
R370 common_bottom.t33 common_bottom.t2 1.2245
R371 common_bottom.t2 common_bottom.t60 1.2245
R372 common_bottom.t51 common_bottom.t60 1.2245
R373 common_bottom.t34 common_bottom.t49 1.2245
R374 common_bottom.t49 common_bottom.t60 1.2245
R375 common_bottom.t49 common_bottom.t19 1.2245
R376 common_bottom.t19 common_bottom.t2 1.2245
R377 common_bottom.t19 common_bottom.t46 1.2245
R378 common_bottom.t46 common_bottom.t33 1.2245
R379 common_bottom.t46 common_bottom.t31 1.2245
R380 common_bottom.t31 common_bottom.t11 1.2245
R381 common_bottom.t16 common_bottom.t3 1.2245
R382 common_bottom.t31 common_bottom.t16 1.2245
R383 common_bottom.t16 common_bottom.t57 1.2245
R384 common_bottom.t8 common_bottom.t43 1.2245
R385 common_bottom.t16 common_bottom.t8 1.2245
R386 common_bottom.t8 common_bottom.t7 1.2245
R387 common_bottom.t48 common_bottom.t32 1.2245
R388 common_bottom.t48 common_bottom.t3 1.2245
R389 common_bottom.t0 common_bottom.t54 1.2245
R390 common_bottom.t0 common_bottom.t13 1.2245
R391 common_bottom.t13 common_bottom.t3 1.2245
R392 common_bottom.t13 common_bottom.t38 1.2245
R393 common_bottom.t38 common_bottom.t14 1.2245
R394 common_bottom.t38 common_bottom.t18 1.2245
R395 common_bottom.t18 common_bottom.t61 1.2245
R396 common_bottom.t18 common_bottom.t12 1.2245
R397 common_bottom.t18 common_bottom.t63 1.2245
R398 common_bottom.t63 common_bottom.t21 1.2245
R399 common_bottom.t63 common_bottom.t24 1.2245
R400 common_bottom.t24 common_bottom.t20 1.2245
R401 common_bottom.t24 common_bottom.t41 1.2245
R402 common_bottom.t41 common_bottom.t55 1.2245
R403 common_bottom.t52 common_bottom.t36 1.2245
R404 common_bottom.t39 common_bottom.t25 1.2245
R405 common_bottom.t24 common_bottom.t25 1.2245
R406 common_bottom.t5 common_bottom.t61 1.2245
R407 common_bottom.t25 common_bottom.t5 1.2245
R408 common_bottom.t63 common_bottom.t5 1.2245
R409 common_bottom.t36 common_bottom.t50 1.2245
R410 common_bottom.t50 common_bottom.t58 1.2245
R411 common_bottom.t47 common_bottom.t22 1.2245
R412 common_bottom.t58 common_bottom.t47 1.2245
R413 common_bottom.t61 common_bottom.t37 1.2245
R414 common_bottom.t38 common_bottom.t37 1.2245
R415 common_bottom.t37 common_bottom.t53 1.2245
R416 common_bottom.t13 common_bottom.t53 1.2245
R417 common_bottom.t1 common_bottom.t35 1.2245
R418 common_bottom.t53 common_bottom.t35 1.2245
R419 common_bottom.t0 common_bottom.t35 1.2245
R420 common_bottom.t22 common_bottom.t9 1.2245
R421 common_bottom.t9 common_bottom.t6 1.2245
R422 common_bottom.t40 common_bottom.t56 1.2245
R423 common_bottom.t28 common_bottom.t40 1.2245
R424 common_bottom.t40 common_bottom.t26 1.2245
R425 common_bottom.t26 common_bottom.t62 1.2245
R426 common_bottom.t26 common_bottom.t23 1.2245
R427 common_bottom.t23 common_bottom.t10 1.2245
R428 common_bottom.t23 common_bottom.t27 1.2245
R429 common_bottom.t27 common_bottom.t44 1.2245
R430 common_bottom.t27 common_bottom.t59 1.2245
R431 common_bottom.t59 common_bottom.t30 1.2245
R432 common_bottom.t59 common_bottom.t4 1.2245
R433 common_bottom.t45 common_bottom.t4 1.2245
R434 common_bottom.t15 common_bottom.t4 1.2245
R435 common_bottom.t15 common_bottom.t17 1.2245
R436 top_c3.n78 top_c3.n77 16.6385
R437 top_c3.n55 top_c3.n54 5.10563
R438 top_c3.n63 top_c3.n62 5.10563
R439 top_c3.n70 top_c3.n69 5.10563
R440 top_c3.n16 top_c3.n15 5.10563
R441 top_c3.n24 top_c3.n23 5.10563
R442 top_c3.n31 top_c3.n30 5.10563
R443 top_c3.n53 top_c3.n50 4.5005
R444 top_c3.n54 top_c3.n53 4.5005
R445 top_c3.n57 top_c3.n55 4.5005
R446 top_c3.n57 top_c3.n56 4.5005
R447 top_c3.n61 top_c3.n47 4.5005
R448 top_c3.n62 top_c3.n61 4.5005
R449 top_c3.n63 top_c3.n44 4.5005
R450 top_c3.n45 top_c3.n44 4.5005
R451 top_c3.n68 top_c3.n43 4.5005
R452 top_c3.n69 top_c3.n68 4.5005
R453 top_c3.n72 top_c3.n70 4.5005
R454 top_c3.n72 top_c3.n71 4.5005
R455 top_c3.n76 top_c3.n40 4.5005
R456 top_c3.n77 top_c3.n76 4.5005
R457 top_c3.n14 top_c3.n11 4.5005
R458 top_c3.n15 top_c3.n14 4.5005
R459 top_c3.n18 top_c3.n16 4.5005
R460 top_c3.n18 top_c3.n17 4.5005
R461 top_c3.n22 top_c3.n8 4.5005
R462 top_c3.n23 top_c3.n22 4.5005
R463 top_c3.n24 top_c3.n5 4.5005
R464 top_c3.n6 top_c3.n5 4.5005
R465 top_c3.n29 top_c3.n4 4.5005
R466 top_c3.n30 top_c3.n29 4.5005
R467 top_c3.n33 top_c3.n31 4.5005
R468 top_c3.n33 top_c3.n32 4.5005
R469 top_c3.n37 top_c3.n1 4.5005
R470 top_c3.n38 top_c3.n37 4.5005
R471 top_c3.n78 top_c3.n38 4.43436
R472 top_c3.n51 top_c3.n50 3.87383
R473 top_c3.n12 top_c3.n11 3.86303
R474 top_c3.n73 top_c3.n41 2.26321
R475 top_c3.n58 top_c3.n48 2.26321
R476 top_c3.n52 top_c3.n49 2.26321
R477 top_c3.n67 top_c3.n42 2.26321
R478 top_c3.n34 top_c3.n2 2.26321
R479 top_c3.n19 top_c3.n9 2.26321
R480 top_c3.n13 top_c3.n10 2.26321
R481 top_c3.n28 top_c3.n3 2.26321
R482 top_c3.n60 top_c3.n46 2.26285
R483 top_c3.n65 top_c3.n64 2.26285
R484 top_c3.n75 top_c3.n39 2.26285
R485 top_c3.n21 top_c3.n7 2.26285
R486 top_c3.n26 top_c3.n25 2.26285
R487 top_c3.n36 top_c3.n0 2.26285
R488 top_c3.n21 top_c3.n20 1.68355
R489 top_c3.n20 top_c3.n19 1.68355
R490 top_c3.n36 top_c3.n35 1.68115
R491 top_c3.n35 top_c3.n34 1.68115
R492 top_c3.n75 top_c3.n74 1.67275
R493 top_c3.n74 top_c3.n73 1.67275
R494 top_c3.n60 top_c3.n59 1.67275
R495 top_c3.n59 top_c3.n58 1.67275
R496 top_c3.n67 top_c3.n66 1.44115
R497 top_c3.n66 top_c3.n65 1.44115
R498 top_c3.n52 top_c3.n51 1.44115
R499 top_c3.n28 top_c3.n27 1.43035
R500 top_c3.n27 top_c3.n26 1.43035
R501 top_c3.n13 top_c3.n12 1.43035
R502 top_c3.n56 top_c3.n47 1.28063
R503 top_c3.n45 top_c3.n43 1.28063
R504 top_c3.n71 top_c3.n40 1.28063
R505 top_c3.n17 top_c3.n8 1.28063
R506 top_c3.n6 top_c3.n4 1.28063
R507 top_c3.n32 top_c3.n1 1.28063
R508 top_c3 top_c3.n78 1.08068
R509 top_c3.n74 top_c3.t5 0.122337
R510 top_c3.n66 top_c3.t2 0.122337
R511 top_c3.n59 top_c3.t6 0.122337
R512 top_c3.n51 top_c3.t4 0.122337
R513 top_c3.n35 top_c3.t7 0.122337
R514 top_c3.n27 top_c3.t1 0.122337
R515 top_c3.n20 top_c3.t0 0.122337
R516 top_c3.n12 top_c3.t3 0.122337
R517 top_c3.n54 top_c3.n49 0.0269027
R518 top_c3.n50 top_c3.n49 0.0269027
R519 top_c3.n56 top_c3.n48 0.0269027
R520 top_c3.n55 top_c3.n48 0.0269027
R521 top_c3.n62 top_c3.n46 0.0269027
R522 top_c3.n47 top_c3.n46 0.0269027
R523 top_c3.n64 top_c3.n45 0.0269027
R524 top_c3.n64 top_c3.n63 0.0269027
R525 top_c3.n69 top_c3.n42 0.0269027
R526 top_c3.n43 top_c3.n42 0.0269027
R527 top_c3.n71 top_c3.n41 0.0269027
R528 top_c3.n70 top_c3.n41 0.0269027
R529 top_c3.n77 top_c3.n39 0.0269027
R530 top_c3.n40 top_c3.n39 0.0269027
R531 top_c3.n15 top_c3.n10 0.0269027
R532 top_c3.n11 top_c3.n10 0.0269027
R533 top_c3.n17 top_c3.n9 0.0269027
R534 top_c3.n16 top_c3.n9 0.0269027
R535 top_c3.n23 top_c3.n7 0.0269027
R536 top_c3.n8 top_c3.n7 0.0269027
R537 top_c3.n25 top_c3.n6 0.0269027
R538 top_c3.n25 top_c3.n24 0.0269027
R539 top_c3.n30 top_c3.n3 0.0269027
R540 top_c3.n4 top_c3.n3 0.0269027
R541 top_c3.n32 top_c3.n2 0.0269027
R542 top_c3.n31 top_c3.n2 0.0269027
R543 top_c3.n38 top_c3.n0 0.0269027
R544 top_c3.n1 top_c3.n0 0.0269027
R545 top_c3.n76 top_c3.n75 0.0256609
R546 top_c3.n65 top_c3.n44 0.0256609
R547 top_c3.n61 top_c3.n60 0.0256609
R548 top_c3.n37 top_c3.n36 0.0256609
R549 top_c3.n26 top_c3.n5 0.0256609
R550 top_c3.n22 top_c3.n21 0.0256609
R551 top_c3.n73 top_c3.n72 0.0253044
R552 top_c3.n68 top_c3.n67 0.0253044
R553 top_c3.n58 top_c3.n57 0.0253044
R554 top_c3.n53 top_c3.n52 0.0253044
R555 top_c3.n34 top_c3.n33 0.0253044
R556 top_c3.n29 top_c3.n28 0.0253044
R557 top_c3.n19 top_c3.n18 0.0253044
R558 top_c3.n14 top_c3.n13 0.0253044
R559 top_c4.n115 top_c4.n114 23.6653
R560 top_c4.n115 top_c4.n57 8.09061
R561 top_c4.n38 top_c4.n37 5.1094
R562 top_c4.n85 top_c4.n84 5.10563
R563 top_c4.n75 top_c4.n69 4.5005
R564 top_c4.n76 top_c4.n75 4.5005
R565 top_c4.n79 top_c4.n77 4.5005
R566 top_c4.n79 top_c4.n78 4.5005
R567 top_c4.n83 top_c4.n66 4.5005
R568 top_c4.n84 top_c4.n83 4.5005
R569 top_c4.n103 top_c4.n85 4.5005
R570 top_c4.n103 top_c4.n102 4.5005
R571 top_c4.n101 top_c4.n86 4.5005
R572 top_c4.n99 top_c4.n86 4.5005
R573 top_c4.n98 top_c4.n87 4.5005
R574 top_c4.n96 top_c4.n87 4.5005
R575 top_c4.n95 top_c4.n88 4.5005
R576 top_c4.n93 top_c4.n88 4.5005
R577 top_c4.n92 top_c4.n89 4.5005
R578 top_c4.n90 top_c4.n89 4.5005
R579 top_c4.n113 top_c4.n59 4.5005
R580 top_c4.n114 top_c4.n113 4.5005
R581 top_c4.n27 top_c4.n12 4.5005
R582 top_c4.n25 top_c4.n12 4.5005
R583 top_c4.n24 top_c4.n13 4.5005
R584 top_c4.n22 top_c4.n13 4.5005
R585 top_c4.n21 top_c4.n14 4.5005
R586 top_c4.n19 top_c4.n14 4.5005
R587 top_c4.n18 top_c4.n15 4.5005
R588 top_c4.n16 top_c4.n15 4.5005
R589 top_c4.n36 top_c4.n7 4.5005
R590 top_c4.n37 top_c4.n36 4.5005
R591 top_c4.n38 top_c4.n5 4.5005
R592 top_c4.n41 top_c4.n38 4.5005
R593 top_c4.n45 top_c4.n4 4.5005
R594 top_c4.n46 top_c4.n45 4.5005
R595 top_c4.n49 top_c4.n47 4.5005
R596 top_c4.n49 top_c4.n48 4.5005
R597 top_c4.n56 top_c4.n1 4.5005
R598 top_c4.n57 top_c4.n56 4.5005
R599 top_c4.n28 top_c4.n27 3.89131
R600 top_c4.n73 top_c4.n69 3.87503
R601 top_c4.n42 top_c4.n41 2.2874
R602 top_c4.n26 top_c4.n11 2.26514
R603 top_c4.n23 top_c4.n10 2.26514
R604 top_c4.n20 top_c4.n9 2.26514
R605 top_c4.n17 top_c4.n8 2.26514
R606 top_c4.n35 top_c4.n6 2.26514
R607 top_c4.n44 top_c4.n3 2.26514
R608 top_c4.n104 top_c4.n64 2.26321
R609 top_c4.n80 top_c4.n67 2.26321
R610 top_c4.n74 top_c4.n68 2.26321
R611 top_c4.n50 top_c4.n2 2.26321
R612 top_c4.n82 top_c4.n65 2.26285
R613 top_c4.n100 top_c4.n63 2.26285
R614 top_c4.n97 top_c4.n62 2.26285
R615 top_c4.n94 top_c4.n61 2.26285
R616 top_c4.n91 top_c4.n60 2.26285
R617 top_c4.n112 top_c4.n58 2.26285
R618 top_c4.n55 top_c4.n0 2.26285
R619 top_c4.n42 top_c4.n5 2.251
R620 top_c4.n40 top_c4.n39 2.23805
R621 top_c4.n47 top_c4.n46 1.73939
R622 top_c4.n25 top_c4.n24 1.73714
R623 top_c4.n19 top_c4.n18 1.73714
R624 top_c4.n77 top_c4.n76 1.73063
R625 top_c4.n99 top_c4.n98 1.73063
R626 top_c4.n93 top_c4.n92 1.73063
R627 top_c4.n105 top_c4.n104 1.70061
R628 top_c4.n82 top_c4.n81 1.70061
R629 top_c4.n81 top_c4.n80 1.70061
R630 top_c4.n106 top_c4.n63 1.67275
R631 top_c4.n109 top_c4.n61 1.67275
R632 top_c4.n107 top_c4.n62 1.67275
R633 top_c4.n111 top_c4.n60 1.67275
R634 top_c4.n112 top_c4.n111 1.67275
R635 top_c4.n55 top_c4.n54 1.67275
R636 top_c4.n54 top_c4.n50 1.67275
R637 top_c4.n35 top_c4.n34 1.47908
R638 top_c4.n44 top_c4.n43 1.4788
R639 top_c4.n28 top_c4.n11 1.45122
R640 top_c4.n30 top_c4.n10 1.45122
R641 top_c4.n32 top_c4.n9 1.45122
R642 top_c4.n33 top_c4.n8 1.45122
R643 top_c4.n74 top_c4.n73 1.44235
R644 top_c4.n48 top_c4.n1 1.29188
R645 top_c4.n22 top_c4.n21 1.28714
R646 top_c4.n16 top_c4.n7 1.28714
R647 top_c4.n39 top_c4.n4 1.28489
R648 top_c4.n78 top_c4.n66 1.28063
R649 top_c4.n102 top_c4.n101 1.28063
R650 top_c4.n96 top_c4.n95 1.28063
R651 top_c4.n90 top_c4.n59 1.28063
R652 top_c4 top_c4.n115 0.810684
R653 top_c4.n70 top_c4.t14 0.586765
R654 top_c4.n51 top_c4.t9 0.586765
R655 top_c4.n72 top_c4.n71 0.5405
R656 top_c4.n53 top_c4.n52 0.5405
R657 top_c4.n71 top_c4.n70 0.526689
R658 top_c4.n52 top_c4.n51 0.526689
R659 top_c4.n107 top_c4.n106 0.484786
R660 top_c4.n33 top_c4.n32 0.484786
R661 top_c4.n30 top_c4.n29 0.483143
R662 top_c4.n110 top_c4.n109 0.482942
R663 top_c4.n43 top_c4.n42 0.356001
R664 top_c4.n110 top_c4.t4 0.113497
R665 top_c4.n70 top_c4.t2 0.106765
R666 top_c4.n51 top_c4.t0 0.106765
R667 top_c4.n29 top_c4.t13 0.106765
R668 top_c4.n108 top_c4.t15 0.0923367
R669 top_c4.n105 top_c4.t5 0.0923367
R670 top_c4.n81 top_c4.t6 0.0923367
R671 top_c4.n71 top_c4.t12 0.0923367
R672 top_c4.n72 top_c4.t3 0.0923367
R673 top_c4.n52 top_c4.t7 0.0923367
R674 top_c4.n53 top_c4.t8 0.0923367
R675 top_c4.n43 top_c4.t10 0.0923367
R676 top_c4.n34 top_c4.t11 0.0923367
R677 top_c4.n31 top_c4.t1 0.0923367
R678 top_c4.n39 top_c4.n38 0.0526053
R679 top_c4.n73 top_c4.n72 0.0305
R680 top_c4.n54 top_c4.n53 0.0297722
R681 top_c4.n108 top_c4.n107 0.0283571
R682 top_c4.n109 top_c4.n108 0.0283571
R683 top_c4.n106 top_c4.n105 0.0283571
R684 top_c4.n34 top_c4.n33 0.0283571
R685 top_c4.n31 top_c4.n30 0.0283571
R686 top_c4.n32 top_c4.n31 0.0283571
R687 top_c4.n45 top_c4.n44 0.0269162
R688 top_c4.n12 top_c4.n11 0.0269149
R689 top_c4.n13 top_c4.n10 0.0269149
R690 top_c4.n14 top_c4.n9 0.0269149
R691 top_c4.n15 top_c4.n8 0.0269149
R692 top_c4.n36 top_c4.n35 0.0269149
R693 top_c4.n76 top_c4.n68 0.0269027
R694 top_c4.n69 top_c4.n68 0.0269027
R695 top_c4.n78 top_c4.n67 0.0269027
R696 top_c4.n77 top_c4.n67 0.0269027
R697 top_c4.n84 top_c4.n65 0.0269027
R698 top_c4.n66 top_c4.n65 0.0269027
R699 top_c4.n102 top_c4.n64 0.0269027
R700 top_c4.n85 top_c4.n64 0.0269027
R701 top_c4.n100 top_c4.n99 0.0269027
R702 top_c4.n101 top_c4.n100 0.0269027
R703 top_c4.n97 top_c4.n96 0.0269027
R704 top_c4.n98 top_c4.n97 0.0269027
R705 top_c4.n94 top_c4.n93 0.0269027
R706 top_c4.n95 top_c4.n94 0.0269027
R707 top_c4.n91 top_c4.n90 0.0269027
R708 top_c4.n92 top_c4.n91 0.0269027
R709 top_c4.n114 top_c4.n58 0.0269027
R710 top_c4.n59 top_c4.n58 0.0269027
R711 top_c4.n40 top_c4.n5 0.0269027
R712 top_c4.n26 top_c4.n25 0.0269027
R713 top_c4.n27 top_c4.n26 0.0269027
R714 top_c4.n23 top_c4.n22 0.0269027
R715 top_c4.n24 top_c4.n23 0.0269027
R716 top_c4.n20 top_c4.n19 0.0269027
R717 top_c4.n21 top_c4.n20 0.0269027
R718 top_c4.n17 top_c4.n16 0.0269027
R719 top_c4.n18 top_c4.n17 0.0269027
R720 top_c4.n37 top_c4.n6 0.0269027
R721 top_c4.n7 top_c4.n6 0.0269027
R722 top_c4.n41 top_c4.n40 0.0269027
R723 top_c4.n46 top_c4.n3 0.0269027
R724 top_c4.n4 top_c4.n3 0.0269027
R725 top_c4.n48 top_c4.n2 0.0269027
R726 top_c4.n47 top_c4.n2 0.0269027
R727 top_c4.n57 top_c4.n0 0.0269027
R728 top_c4.n1 top_c4.n0 0.0269027
R729 top_c4.n86 top_c4.n63 0.0256609
R730 top_c4.n88 top_c4.n61 0.0256609
R731 top_c4.n87 top_c4.n62 0.0256609
R732 top_c4.n89 top_c4.n60 0.0256609
R733 top_c4.n113 top_c4.n112 0.0256609
R734 top_c4.n83 top_c4.n82 0.0256609
R735 top_c4.n56 top_c4.n55 0.0256609
R736 top_c4.n104 top_c4.n103 0.0253044
R737 top_c4.n80 top_c4.n79 0.0253044
R738 top_c4.n75 top_c4.n74 0.0253044
R739 top_c4.n50 top_c4.n49 0.0253044
R740 top_c4.n111 top_c4.n110 0.0171124
R741 top_c4.n29 top_c4.n28 0.0166786
R742 top_c0 top_c0.n16 15.7278
R743 top_c0.n8 top_c0.n5 4.5005
R744 top_c0.n9 top_c0.n8 4.5005
R745 top_c0.n10 top_c0.n2 4.5005
R746 top_c0.n3 top_c0.n2 4.5005
R747 top_c0.n15 top_c0.n1 4.5005
R748 top_c0.n16 top_c0.n15 4.5005
R749 top_c0.n6 top_c0.n5 3.86303
R750 top_c0.n7 top_c0.n4 2.26321
R751 top_c0.n14 top_c0.n0 2.26321
R752 top_c0.n12 top_c0.n11 2.26285
R753 top_c0.n10 top_c0.n9 1.73063
R754 top_c0.n14 top_c0.n13 1.43035
R755 top_c0.n13 top_c0.n12 1.43035
R756 top_c0.n7 top_c0.n6 1.43035
R757 top_c0.n3 top_c0.n1 1.28063
R758 top_c0.n13 top_c0.t0 0.122337
R759 top_c0.n6 top_c0.t1 0.122337
R760 top_c0.n9 top_c0.n4 0.0269027
R761 top_c0.n5 top_c0.n4 0.0269027
R762 top_c0.n11 top_c0.n3 0.0269027
R763 top_c0.n11 top_c0.n10 0.0269027
R764 top_c0.n16 top_c0.n0 0.0269027
R765 top_c0.n1 top_c0.n0 0.0269027
R766 top_c0.n12 top_c0.n2 0.0256609
R767 top_c0.n15 top_c0.n14 0.0253044
R768 top_c0.n8 top_c0.n7 0.0253044
R769 top_c2.n20 top_c2.t0 13.6405
R770 top_c2.n28 top_c2.n27 13.5077
R771 top_c2.n28 top_c2.n16 10.8694
R772 top_c2.n10 top_c2.n9 8.48063
R773 top_c2.n22 top_c2.n20 4.5005
R774 top_c2.n22 top_c2.n21 4.5005
R775 top_c2.n26 top_c2.n18 4.5005
R776 top_c2.n27 top_c2.n26 4.5005
R777 top_c2.n8 top_c2.n5 4.5005
R778 top_c2.n9 top_c2.n8 4.5005
R779 top_c2.n10 top_c2.n2 4.5005
R780 top_c2.n3 top_c2.n2 4.5005
R781 top_c2.n15 top_c2.n1 4.5005
R782 top_c2.n16 top_c2.n15 4.5005
R783 top_c2.n6 top_c2.n5 3.86303
R784 top_c2.n23 top_c2.n19 2.26321
R785 top_c2.n7 top_c2.n4 2.26321
R786 top_c2.n14 top_c2.n0 2.26321
R787 top_c2.n25 top_c2.n17 2.26285
R788 top_c2.n12 top_c2.n11 2.26285
R789 top_c2.n14 top_c2.n13 1.43035
R790 top_c2.n13 top_c2.n12 1.43035
R791 top_c2.n7 top_c2.n6 1.43035
R792 top_c2.n25 top_c2.n24 1.37695
R793 top_c2.n24 top_c2.n23 1.37695
R794 top_c2 top_c2.n28 1.37431
R795 top_c2.n21 top_c2.n18 1.28063
R796 top_c2.n3 top_c2.n1 1.28063
R797 top_c2.n24 top_c2.t2 0.122337
R798 top_c2.n13 top_c2.t3 0.122337
R799 top_c2.n6 top_c2.t1 0.122337
R800 top_c2.n21 top_c2.n19 0.0269027
R801 top_c2.n20 top_c2.n19 0.0269027
R802 top_c2.n27 top_c2.n17 0.0269027
R803 top_c2.n18 top_c2.n17 0.0269027
R804 top_c2.n9 top_c2.n4 0.0269027
R805 top_c2.n5 top_c2.n4 0.0269027
R806 top_c2.n11 top_c2.n3 0.0269027
R807 top_c2.n11 top_c2.n10 0.0269027
R808 top_c2.n16 top_c2.n0 0.0269027
R809 top_c2.n1 top_c2.n0 0.0269027
R810 top_c2.n26 top_c2.n25 0.0256609
R811 top_c2.n12 top_c2.n2 0.0256609
R812 top_c2.n23 top_c2.n22 0.0253044
R813 top_c2.n15 top_c2.n14 0.0253044
R814 top_c2.n8 top_c2.n7 0.0253044
R815 top_c_dummy top_c_dummy.n5 12.3767
R816 top_c_dummy.n4 top_c_dummy.n1 4.5005
R817 top_c_dummy.n5 top_c_dummy.n4 4.5005
R818 top_c_dummy.n2 top_c_dummy.n1 3.87863
R819 top_c_dummy.n3 top_c_dummy.n0 2.26285
R820 top_c_dummy.n3 top_c_dummy.n2 1.44595
R821 top_c_dummy.n2 top_c_dummy.t0 0.122337
R822 top_c_dummy.n5 top_c_dummy.n0 0.0269027
R823 top_c_dummy.n1 top_c_dummy.n0 0.0269027
R824 top_c_dummy.n4 top_c_dummy.n3 0.0256609
R825 top_c1 top_c1.n5 8.97918
R826 top_c1.n4 top_c1.n1 4.5005
R827 top_c1.n5 top_c1.n4 4.5005
R828 top_c1.n2 top_c1.n1 3.80963
R829 top_c1.n3 top_c1.n0 2.26285
R830 top_c1.n3 top_c1.n2 1.37695
R831 top_c1.n2 top_c1.t0 0.122337
R832 top_c1.n5 top_c1.n0 0.0269027
R833 top_c1.n1 top_c1.n0 0.0269027
R834 top_c1.n4 top_c1.n3 0.0256609
C0 top_c3 common_bottom 11.1152f
C1 common_bottom m3_1090_37400 0.97368f
C2 top_c5 top_c2 2.34498f
C3 top_c1 top_c4 0.47261f
C4 top_c5 common_bottom 33.806698f
C5 m3_16090_37400 common_bottom 0.971673f
C6 top_c3 top_c0 0.200626f
C7 m3_9610_37600 top_c2 3.19116f
C8 top_c5 top_c0 0.971104f
C9 common_bottom m3_9610_37600 0.97376f
C10 top_c_dummy top_c1 0.013558f
C11 top_c3 m3_1090_37400 3.45276f
C12 m3_n1905_37400 top_c4 3.43141f
C13 top_c_dummy top_c4 0.491368f
C14 top_c3 top_c5 3.3804f
C15 top_c3 m3_16090_37400 0.017098f
C16 top_c5 m3_1090_37400 0.432815f
C17 top_c5 m3_16090_37400 0.590451f
C18 m3_13080_37400 top_c4 0.177159f
C19 top_c3 m3_9610_37600 0.026795f
C20 top_c1 top_c2 0.077876f
C21 common_bottom top_c1 2.13473f
C22 top_c5 m3_9610_37600 0.683089f
C23 top_c2 top_c4 0.741784f
C24 common_bottom top_c4 18.375599f
C25 top_c1 top_c0 3.33484f
C26 top_c_dummy top_c2 3.76834f
C27 top_c0 top_c4 0.520991f
C28 m3_n1905_37400 common_bottom 0.977097f
C29 top_c3 top_c1 0.200621f
C30 common_bottom top_c_dummy 2.08325f
C31 top_c3 top_c4 5.20067f
C32 m3_1090_37400 top_c4 0.152828f
C33 top_c5 top_c1 1.05695f
C34 m3_13080_37400 top_c2 0.028837f
C35 top_c5 top_c4 9.36867f
C36 m3_16090_37400 top_c4 3.84867f
C37 common_bottom m3_13080_37400 1.11039f
C38 top_c_dummy top_c0 0.569f
C39 top_c3 m3_n1905_37400 0.245343f
C40 top_c1 m3_9610_37600 0.135476f
C41 top_c3 top_c_dummy 0.084329f
C42 common_bottom top_c2 6.94043f
C43 m3_9610_37600 top_c4 0.290507f
C44 top_c5 m3_n1905_37400 0.719426f
C45 top_c5 top_c_dummy 0.619868f
C46 top_c3 m3_13080_37400 3.66429f
C47 top_c0 top_c2 0.090243f
C48 common_bottom top_c0 3.29289f
C49 top_c5 m3_13080_37400 0.804262f
C50 top_c3 top_c2 3.15711f
C51 m3_1090_37400 top_c2 0.27095f
C52 common_bottom VSUBS 80.35331f
C53 top_c1 VSUBS 7.865008f
C54 top_c0 VSUBS 9.978719f
C55 top_c_dummy VSUBS 8.040878f
C56 top_c2 VSUBS 19.660772f
C57 top_c3 VSUBS 29.157608f
C58 top_c5 VSUBS 85.81033f
C59 top_c4 VSUBS 45.84397f
C60 m3_16090_37400 VSUBS 4.73364f $ **FLOATING
C61 m3_13080_37400 VSUBS 4.84066f $ **FLOATING
C62 m3_9610_37600 VSUBS 4.70657f $ **FLOATING
C63 m3_1090_37400 VSUBS 4.77027f $ **FLOATING
C64 m3_n1905_37400 VSUBS 4.74427f $ **FLOATING
C65 top_c1.n1 VSUBS -1.04934f
C66 top_c1.t0 VSUBS 3.63772f
C67 top_c1.n2 VSUBS 1.65722f
C68 top_c1.n3 VSUBS 0.047436f
C69 top_c1.n4 VSUBS 0.031183f
C70 top_c1.n5 VSUBS 0.546014f
C71 top_c_dummy.n1 VSUBS -0.759566f
C72 top_c_dummy.t0 VSUBS 3.45403f
C73 top_c_dummy.n2 VSUBS 1.73536f
C74 top_c_dummy.n3 VSUBS 0.050426f
C75 top_c_dummy.n4 VSUBS 0.029608f
C76 top_c_dummy.n5 VSUBS 0.704013f
C77 top_c2.n1 VSUBS 0.069098f
C78 top_c2.t3 VSUBS 2.4961f
C79 top_c2.n2 VSUBS 0.021397f
C80 top_c2.n3 VSUBS 0.070776f
C81 top_c2.n5 VSUBS -0.019384f
C82 top_c2.t1 VSUBS 2.4961f
C83 top_c2.n6 VSUBS 1.51897f
C84 top_c2.n7 VSUBS 0.035839f
C85 top_c2.n8 VSUBS 0.021092f
C86 top_c2.n9 VSUBS 0.354989f
C87 top_c2.n10 VSUBS 0.353262f
C88 top_c2.n12 VSUBS 0.03554f
C89 top_c2.n13 VSUBS 1.54005f
C90 top_c2.n14 VSUBS 0.035839f
C91 top_c2.n15 VSUBS 0.021092f
C92 top_c2.n16 VSUBS 0.449324f
C93 top_c2.n18 VSUBS 0.069098f
C94 top_c2.t2 VSUBS 2.4961f
C95 top_c2.t0 VSUBS 3.84401f
C96 top_c2.n20 VSUBS 0.279175f
C97 top_c2.n21 VSUBS 0.070776f
C98 top_c2.n22 VSUBS 0.021092f
C99 top_c2.n23 VSUBS 0.032848f
C100 top_c2.n24 VSUBS 1.52627f
C101 top_c2.n25 VSUBS 0.032549f
C102 top_c2.n26 VSUBS 0.021397f
C103 top_c2.n27 VSUBS 0.472165f
C104 top_c2.n28 VSUBS 0.97149f
C105 top_c0.n1 VSUBS 0.047889f
C106 top_c0.t0 VSUBS 1.72993f
C107 top_c0.n2 VSUBS 0.014829f
C108 top_c0.n3 VSUBS 0.049051f
C109 top_c0.n5 VSUBS -0.135571f
C110 top_c0.t1 VSUBS 1.72993f
C111 top_c0.n6 VSUBS 0.990212f
C112 top_c0.n7 VSUBS 0.024838f
C113 top_c0.n8 VSUBS 0.014618f
C114 top_c0.n9 VSUBS 0.061366f
C115 top_c0.n10 VSUBS 0.060193f
C116 top_c0.n12 VSUBS 0.024631f
C117 top_c0.n13 VSUBS 1.06733f
C118 top_c0.n14 VSUBS 0.024838f
C119 top_c0.n15 VSUBS 0.014618f
C120 top_c0.n16 VSUBS 0.444289f
C121 top_c4.n1 VSUBS 0.035791f
C122 top_c4.n4 VSUBS 0.035634f
C123 top_c4.n5 VSUBS 0.010341f
C124 top_c4.n7 VSUBS 0.03568f
C125 top_c4.n8 VSUBS 0.018196f
C126 top_c4.n9 VSUBS 0.018196f
C127 top_c4.n10 VSUBS 0.018196f
C128 top_c4.t13 VSUBS 1.23602f
C129 top_c4.n11 VSUBS 0.018196f
C130 top_c4.n12 VSUBS 0.010341f
C131 top_c4.n13 VSUBS 0.010341f
C132 top_c4.n14 VSUBS 0.010341f
C133 top_c4.n15 VSUBS 0.010341f
C134 top_c4.n16 VSUBS 0.03568f
C135 top_c4.n18 VSUBS 0.044821f
C136 top_c4.n19 VSUBS 0.044821f
C137 top_c4.n21 VSUBS 0.03568f
C138 top_c4.n22 VSUBS 0.03568f
C139 top_c4.n24 VSUBS 0.044821f
C140 top_c4.n25 VSUBS 0.044821f
C141 top_c4.n27 VSUBS 0.077149f
C142 top_c4.n28 VSUBS 0.420531f
C143 top_c4.n29 VSUBS 0.783293f
C144 top_c4.n30 VSUBS 0.442984f
C145 top_c4.t1 VSUBS 1.11982f
C146 top_c4.n31 VSUBS 0.519914f
C147 top_c4.n32 VSUBS 0.433775f
C148 top_c4.n33 VSUBS 0.433775f
C149 top_c4.t11 VSUBS 1.11982f
C150 top_c4.n34 VSUBS 0.775103f
C151 top_c4.n35 VSUBS 0.023097f
C152 top_c4.n36 VSUBS 0.010341f
C153 top_c4.n37 VSUBS 0.113403f
C154 top_c4.n38 VSUBS 0.113473f
C155 top_c4.n39 VSUBS 0.035634f
C156 top_c4.n41 VSUBS 0.010526f
C157 top_c4.n42 VSUBS 0.052632f
C158 top_c4.t10 VSUBS 1.11982f
C159 top_c4.n43 VSUBS 0.990253f
C160 top_c4.n44 VSUBS 0.023088f
C161 top_c4.n45 VSUBS 0.010341f
C162 top_c4.n46 VSUBS 0.044867f
C163 top_c4.n47 VSUBS 0.044867f
C164 top_c4.n48 VSUBS 0.036654f
C165 top_c4.n49 VSUBS 0.010855f
C166 top_c4.n50 VSUBS 0.026238f
C167 top_c4.t0 VSUBS 1.22058f
C168 top_c4.t9 VSUBS 1.92787f
C169 top_c4.n51 VSUBS 1.19931f
C170 top_c4.t7 VSUBS 1.11982f
C171 top_c4.n52 VSUBS 1.13247f
C172 top_c4.t8 VSUBS 1.11982f
C173 top_c4.n53 VSUBS 0.842042f
C174 top_c4.n54 VSUBS 0.401937f
C175 top_c4.n55 VSUBS 0.026085f
C176 top_c4.n56 VSUBS 0.011012f
C177 top_c4.n57 VSUBS 0.174811f
C178 top_c4.n59 VSUBS 0.035562f
C179 top_c4.n60 VSUBS 0.026085f
C180 top_c4.n61 VSUBS 0.026085f
C181 top_c4.n62 VSUBS 0.026085f
C182 top_c4.n63 VSUBS 0.026085f
C183 top_c4.n66 VSUBS 0.035562f
C184 top_c4.n69 VSUBS -0.100752f
C185 top_c4.t2 VSUBS 1.22058f
C186 top_c4.t14 VSUBS 1.92787f
C187 top_c4.n70 VSUBS 1.19931f
C188 top_c4.t12 VSUBS 1.11982f
C189 top_c4.n71 VSUBS 1.13247f
C190 top_c4.t3 VSUBS 1.11982f
C191 top_c4.n72 VSUBS 0.843126f
C192 top_c4.n73 VSUBS 0.232738f
C193 top_c4.n74 VSUBS 0.018801f
C194 top_c4.n75 VSUBS 0.010855f
C195 top_c4.n76 VSUBS 0.045571f
C196 top_c4.n77 VSUBS 0.0447f
C197 top_c4.n78 VSUBS 0.036426f
C198 top_c4.n79 VSUBS 0.010855f
C199 top_c4.n80 VSUBS 0.030747f
C200 top_c4.t6 VSUBS 1.11982f
C201 top_c4.n81 VSUBS 1.06128f
C202 top_c4.n82 VSUBS 0.030594f
C203 top_c4.n83 VSUBS 0.011012f
C204 top_c4.n84 VSUBS 0.114138f
C205 top_c4.n85 VSUBS 0.113253f
C206 top_c4.n86 VSUBS 0.011012f
C207 top_c4.n87 VSUBS 0.011012f
C208 top_c4.n88 VSUBS 0.011012f
C209 top_c4.n89 VSUBS 0.011012f
C210 top_c4.n90 VSUBS 0.036426f
C211 top_c4.n92 VSUBS 0.0447f
C212 top_c4.n93 VSUBS 0.045571f
C213 top_c4.n95 VSUBS 0.035562f
C214 top_c4.n96 VSUBS 0.036426f
C215 top_c4.n98 VSUBS 0.0447f
C216 top_c4.n99 VSUBS 0.045571f
C217 top_c4.n101 VSUBS 0.035562f
C218 top_c4.n102 VSUBS 0.036426f
C219 top_c4.n103 VSUBS 0.010855f
C220 top_c4.n104 VSUBS 0.030747f
C221 top_c4.t5 VSUBS 1.11982f
C222 top_c4.n105 VSUBS 0.790595f
C223 top_c4.n106 VSUBS 0.448875f
C224 top_c4.n107 VSUBS 0.448875f
C225 top_c4.t15 VSUBS 1.11982f
C226 top_c4.n108 VSUBS 0.519914f
C227 top_c4.n109 VSUBS 0.45818f
C228 top_c4.t4 VSUBS 1.19845f
C229 top_c4.n110 VSUBS 0.811033f
C230 top_c4.n111 VSUBS 0.427282f
C231 top_c4.n112 VSUBS 0.026085f
C232 top_c4.n113 VSUBS 0.011012f
C233 top_c4.n114 VSUBS 0.457697f
C234 top_c4.n115 VSUBS 0.654605f
C235 top_c3.n1 VSUBS 0.052838f
C236 top_c3.t7 VSUBS 1.90873f
C237 top_c3.n4 VSUBS 0.052838f
C238 top_c3.t1 VSUBS 1.90873f
C239 top_c3.n5 VSUBS 0.016362f
C240 top_c3.n6 VSUBS 0.054121f
C241 top_c3.n8 VSUBS 0.052838f
C242 top_c3.t0 VSUBS 1.90873f
C243 top_c3.n11 VSUBS 0.115446f
C244 top_c3.t3 VSUBS 1.93012f
C245 top_c3.n12 VSUBS 1.35044f
C246 top_c3.n13 VSUBS 0.027405f
C247 top_c3.n14 VSUBS 0.016129f
C248 top_c3.n15 VSUBS 0.169586f
C249 top_c3.n16 VSUBS 0.16827f
C250 top_c3.n17 VSUBS 0.054121f
C251 top_c3.n18 VSUBS 0.016129f
C252 top_c3.n19 VSUBS 0.039538f
C253 top_c3.n20 VSUBS 1.22503f
C254 top_c3.n21 VSUBS 0.03931f
C255 top_c3.n22 VSUBS 0.016362f
C256 top_c3.n23 VSUBS 0.169586f
C257 top_c3.n24 VSUBS 0.16827f
C258 top_c3.n26 VSUBS 0.027177f
C259 top_c3.n27 VSUBS 1.17765f
C260 top_c3.n28 VSUBS 0.027405f
C261 top_c3.n29 VSUBS 0.016129f
C262 top_c3.n30 VSUBS 0.169586f
C263 top_c3.n31 VSUBS 0.16827f
C264 top_c3.n32 VSUBS 0.054121f
C265 top_c3.n33 VSUBS 0.016129f
C266 top_c3.n34 VSUBS 0.039414f
C267 top_c3.n35 VSUBS 1.2246f
C268 top_c3.n36 VSUBS 0.039186f
C269 top_c3.n37 VSUBS 0.016362f
C270 top_c3.n38 VSUBS 0.149418f
C271 top_c3.n40 VSUBS 0.052838f
C272 top_c3.t5 VSUBS 1.94283f
C273 top_c3.n43 VSUBS 0.052838f
C274 top_c3.t2 VSUBS 1.90873f
C275 top_c3.n44 VSUBS 0.016362f
C276 top_c3.n45 VSUBS 0.054121f
C277 top_c3.n47 VSUBS 0.052838f
C278 top_c3.t6 VSUBS 1.9267f
C279 top_c3.n50 VSUBS -0.014712f
C280 top_c3.t4 VSUBS 1.90873f
C281 top_c3.n51 VSUBS 1.164f
C282 top_c3.n52 VSUBS 0.027881f
C283 top_c3.n53 VSUBS 0.016129f
C284 top_c3.n54 VSUBS 0.169586f
C285 top_c3.n55 VSUBS 0.16827f
C286 top_c3.n56 VSUBS 0.054121f
C287 top_c3.n57 VSUBS 0.016129f
C288 top_c3.n58 VSUBS 0.038984f
C289 top_c3.n59 VSUBS 1.27811f
C290 top_c3.n60 VSUBS 0.038756f
C291 top_c3.n61 VSUBS 0.016362f
C292 top_c3.n62 VSUBS 0.169586f
C293 top_c3.n63 VSUBS 0.16827f
C294 top_c3.n65 VSUBS 0.027653f
C295 top_c3.n66 VSUBS 1.17975f
C296 top_c3.n67 VSUBS 0.027881f
C297 top_c3.n68 VSUBS 0.016129f
C298 top_c3.n69 VSUBS 0.169586f
C299 top_c3.n70 VSUBS 0.16827f
C300 top_c3.n71 VSUBS 0.054121f
C301 top_c3.n72 VSUBS 0.016129f
C302 top_c3.n73 VSUBS 0.038984f
C303 top_c3.n74 VSUBS 1.38422f
C304 top_c3.n75 VSUBS 0.038756f
C305 top_c3.n76 VSUBS 0.016362f
C306 top_c3.n77 VSUBS 0.451776f
C307 top_c3.n78 VSUBS 0.656944f
C308 common_bottom.t4 VSUBS 1.16727f
C309 common_bottom.t45 VSUBS 1.2507f
C310 common_bottom.t60 VSUBS 1.25388f
C311 common_bottom.t55 VSUBS 1.16568f
C312 common_bottom.t20 VSUBS 1.2507f
C313 common_bottom.t21 VSUBS 1.2507f
C314 common_bottom.t2 VSUBS 1.25388f
C315 common_bottom.t12 VSUBS 1.2507f
C316 common_bottom.t33 VSUBS 1.25388f
C317 common_bottom.t14 VSUBS 1.2507f
C318 common_bottom.t11 VSUBS 1.25388f
C319 common_bottom.t3 VSUBS 1.25229f
C320 common_bottom.t57 VSUBS 1.25388f
C321 common_bottom.t43 VSUBS 1.16727f
C322 common_bottom.t29 VSUBS 1.16727f
C323 common_bottom.t62 VSUBS 1.2507f
C324 common_bottom.t42 VSUBS 1.16568f
C325 common_bottom.t56 VSUBS 1.08384f
C326 common_bottom.t10 VSUBS 1.2507f
C327 common_bottom.t44 VSUBS 1.2507f
C328 common_bottom.t30 VSUBS 1.2507f
C329 common_bottom.t59 VSUBS 1.16727f
C330 common_bottom.t27 VSUBS 1.16727f
C331 common_bottom.t23 VSUBS 1.16727f
C332 common_bottom.t26 VSUBS 1.16727f
C333 common_bottom.t40 VSUBS 1.16727f
C334 common_bottom.t28 VSUBS 1.2507f
C335 common_bottom.t7 VSUBS 1.25388f
C336 common_bottom.t32 VSUBS 1.16727f
C337 common_bottom.t54 VSUBS 1.16727f
C338 common_bottom.t35 VSUBS 1.2507f
C339 common_bottom.t53 VSUBS 1.25388f
C340 common_bottom.t37 VSUBS 1.25388f
C341 common_bottom.t61 VSUBS 1.2507f
C342 common_bottom.t5 VSUBS 1.2507f
C343 common_bottom.t25 VSUBS 1.25388f
C344 common_bottom.t1 VSUBS 1.16727f
C345 common_bottom.t6 VSUBS 1.08225f
C346 common_bottom.t9 VSUBS 1.16886f
C347 common_bottom.t22 VSUBS 1.16568f
C348 common_bottom.t47 VSUBS 1.16568f
C349 common_bottom.t58 VSUBS 1.16886f
C350 common_bottom.t50 VSUBS 1.16886f
C351 common_bottom.t36 VSUBS 1.16568f
C352 common_bottom.t52 VSUBS 1.08066f
C353 common_bottom.t39 VSUBS 1.17045f
C354 common_bottom.t41 VSUBS 1.16568f
C355 common_bottom.t24 VSUBS 1.25229f
C356 common_bottom.t63 VSUBS 1.25229f
C357 common_bottom.t18 VSUBS 1.25229f
C358 common_bottom.t38 VSUBS 1.25229f
C359 common_bottom.t13 VSUBS 1.25229f
C360 common_bottom.t0 VSUBS 1.25388f
C361 common_bottom.t48 VSUBS 1.25229f
C362 common_bottom.t8 VSUBS 1.2507f
C363 common_bottom.t16 VSUBS 1.25229f
C364 common_bottom.t31 VSUBS 1.25388f
C365 common_bottom.t46 VSUBS 1.25388f
C366 common_bottom.t19 VSUBS 1.25388f
C367 common_bottom.t49 VSUBS 1.25388f
C368 common_bottom.t34 VSUBS 1.17045f
C369 common_bottom.t51 VSUBS 1.16727f
C370 common_bottom.t17 VSUBS 1.16568f
C371 common_bottom.t15 VSUBS 1.21451f
C372 top_c5.n2 VSUBS 0.075379f
C373 top_c5.n9 VSUBS 0.075379f
C374 top_c5.t6 VSUBS 0.692975f
C375 top_c5.n16 VSUBS 0.487389f
C376 top_c5.n17 VSUBS 0.201528f
C377 top_c5.t31 VSUBS 0.692975f
C378 top_c5.n18 VSUBS 0.618598f
C379 top_c5.t7 VSUBS 0.692975f
C380 top_c5.n19 VSUBS 0.58905f
C381 top_c5.t5 VSUBS 1.25799f
C382 top_c5.n20 VSUBS 0.387458f
C383 top_c5.t22 VSUBS 0.692975f
C384 top_c5.n21 VSUBS 0.321738f
C385 top_c5.n22 VSUBS 0.286139f
C386 top_c5.t1 VSUBS 0.692975f
C387 top_c5.n23 VSUBS 0.743412f
C388 top_c5.t15 VSUBS 0.692975f
C389 top_c5.n24 VSUBS 0.743412f
C390 top_c5.n25 VSUBS 0.286997f
C391 top_c5.t17 VSUBS 0.692975f
C392 top_c5.n26 VSUBS 0.321738f
C393 top_c5.n27 VSUBS 0.274351f
C394 top_c5.t4 VSUBS 0.692975f
C395 top_c5.n28 VSUBS 0.321738f
C396 top_c5.n29 VSUBS 0.270472f
C397 top_c5.n30 VSUBS 0.196011f
C398 top_c5.t20 VSUBS 0.692975f
C399 top_c5.n31 VSUBS 0.321738f
C400 top_c5.n32 VSUBS 0.229795f
C401 top_c5.n33 VSUBS 0.249023f
C402 top_c5.n39 VSUBS 0.204314f
C403 top_c5.t21 VSUBS 0.692975f
C404 top_c5.n40 VSUBS 0.597708f
C405 top_c5.t3 VSUBS 0.692975f
C406 top_c5.n41 VSUBS 0.321738f
C407 top_c5.n42 VSUBS 0.22556f
C408 top_c5.t18 VSUBS 1.19021f
C409 top_c5.n43 VSUBS 0.344584f
C410 top_c5.t19 VSUBS 0.692975f
C411 top_c5.n44 VSUBS 0.321738f
C412 top_c5.n45 VSUBS 0.25542f
C413 top_c5.t9 VSUBS 0.692975f
C414 top_c5.n46 VSUBS 0.511347f
C415 top_c5.n47 VSUBS 0.309932f
C416 top_c5.n49 VSUBS 0.213754f
C417 top_c5.n53 VSUBS 0.037725f
C418 top_c5.n55 VSUBS 0.067883f
C419 top_c5.n56 VSUBS 0.067925f
C420 top_c5.n60 VSUBS 0.037725f
C421 top_c5.n62 VSUBS 0.010238f
C422 top_c5.n63 VSUBS 0.010197f
C423 top_c5.n67 VSUBS 0.037725f
C424 top_c5.n69 VSUBS 0.025442f
C425 top_c5.n70 VSUBS 0.025442f
C426 top_c5.n74 VSUBS 0.037725f
C427 top_c5.n76 VSUBS 0.010182f
C428 top_c5.n77 VSUBS 0.010182f
C429 top_c5.n81 VSUBS 0.037725f
C430 top_c5.n83 VSUBS 0.025456f
C431 top_c5.n84 VSUBS 0.025456f
C432 top_c5.n88 VSUBS 0.037725f
C433 top_c5.n90 VSUBS 0.010182f
C434 top_c5.n91 VSUBS 0.010182f
C435 top_c5.n95 VSUBS 0.037725f
C436 top_c5.n97 VSUBS 0.023041f
C437 top_c5.n102 VSUBS 0.226417f
C438 top_c5.t11 VSUBS 0.692975f
C439 top_c5.n103 VSUBS 0.717552f
C440 top_c5.t26 VSUBS 0.692975f
C441 top_c5.n104 VSUBS 0.321738f
C442 top_c5.n105 VSUBS 0.198025f
C443 top_c5.t10 VSUBS 0.755334f
C444 top_c5.t25 VSUBS 1.19302f
C445 top_c5.n106 VSUBS 0.74217f
C446 top_c5.t23 VSUBS 0.692975f
C447 top_c5.n107 VSUBS 0.690402f
C448 top_c5.n108 VSUBS 0.25542f
C449 top_c5.t12 VSUBS 0.692975f
C450 top_c5.n109 VSUBS 0.321738f
C451 top_c5.n110 VSUBS 0.25542f
C452 top_c5.t29 VSUBS 0.692975f
C453 top_c5.n111 VSUBS 0.511347f
C454 top_c5.n117 VSUBS 0.037725f
C455 top_c5.n118 VSUBS 0.305192f
C456 top_c5.n119 VSUBS 0.037725f
C457 top_c5.n123 VSUBS 0.037725f
C458 top_c5.n126 VSUBS 0.037725f
C459 top_c5.n132 VSUBS 0.010182f
C460 top_c5.n133 VSUBS 0.010182f
C461 top_c5.n139 VSUBS 0.025456f
C462 top_c5.n140 VSUBS 0.025456f
C463 top_c5.n146 VSUBS 0.010197f
C464 top_c5.n147 VSUBS 0.010197f
C465 top_c5.n153 VSUBS 0.025442f
C466 top_c5.n154 VSUBS 0.025442f
C467 top_c5.n160 VSUBS 0.030626f
C468 top_c5.n161 VSUBS 0.124905f
C469 top_c5.n162 VSUBS 0.201528f
C470 top_c5.t0 VSUBS 0.692975f
C471 top_c5.n163 VSUBS 0.321738f
C472 top_c5.t28 VSUBS 0.692975f
C473 top_c5.n164 VSUBS 0.737409f
C474 top_c5.t8 VSUBS 0.692975f
C475 top_c5.n165 VSUBS 0.58905f
C476 top_c5.t2 VSUBS 1.31855f
C477 top_c5.n166 VSUBS 0.398317f
C478 top_c5.t24 VSUBS 0.692975f
C479 top_c5.n167 VSUBS 0.321738f
C480 top_c5.n168 VSUBS 0.286139f
C481 top_c5.t13 VSUBS 0.692975f
C482 top_c5.n169 VSUBS 0.743412f
C483 top_c5.t27 VSUBS 0.692975f
C484 top_c5.n170 VSUBS 0.743412f
C485 top_c5.n171 VSUBS 0.286139f
C486 top_c5.t14 VSUBS 0.692975f
C487 top_c5.n172 VSUBS 0.321738f
C488 top_c5.n173 VSUBS 0.278729f
C489 top_c5.n174 VSUBS 0.270541f
C490 top_c5.t16 VSUBS 0.692975f
C491 top_c5.n175 VSUBS 0.326954f
C492 top_c5.n176 VSUBS 0.291674f
C493 top_c5.t30 VSUBS 0.692975f
C494 top_c5.n177 VSUBS 0.455414f
C495 top_c5.n178 VSUBS 0.176072f
C496 top_c5.n179 VSUBS 0.075379f
C497 top_c5.n180 VSUBS 0.037725f
C498 top_c5.n182 VSUBS 0.067883f
C499 top_c5.n183 VSUBS 0.067925f
C500 top_c5.n187 VSUBS 0.010182f
C501 top_c5.n188 VSUBS 0.010224f
C502 top_c5.n193 VSUBS 0.037725f
C503 top_c5.n194 VSUBS 0.188972f
C504 top_c5.n195 VSUBS 0.037725f
C505 top_c5.n197 VSUBS 0.501567f
C506 top_c5.n198 VSUBS 0.524685f
.ends

