* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt TOP S R GND VDD Qn Q
X0 Q.t2 Qn.t3 GND.t3 GND.t2 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X1 GND.t5 S.t0 Qn.t0 GND.t4 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X2 Q.t0 R.t0 GND.t1 GND.t0 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X3 VDD.t3 Q.t3 Qn.t1 VDD.t2 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
X4 GND.t7 Q.t4 Qn.t2 GND.t6 nfet_03v3 ad=1.708p pd=6.82u as=1.708p ps=6.82u w=2.8u l=0.28u
X5 Q.t1 Qn.t4 VDD.t1 VDD.t0 pfet_03v3 ad=1.82p pd=6.9u as=1.82p ps=6.9u w=2.8u l=0.28u
R0 Qn Qn.t4 56.0856
R1 Qn.n1 Qn.t3 55.9719
R2 Qn.n2 Qn.t0 4.35469
R3 Qn.n1 Qn.n0 3.18045
R4 Qn.n0 Qn.t1 3.0207
R5 Qn.n0 Qn.t2 2.1605
R6 Qn.n2 Qn.n1 0.068
R7 Qn Qn.n2 0.0573421
R8 GND.n4 GND.n3 31769.5
R9 GND.n3 GND.n2 31754.7
R10 GND.n9 GND.n3 9378.27
R11 GND.n9 GND.t6 1534.44
R12 GND.t2 GND.n9 1534.44
R13 GND.t6 GND.n8 854.365
R14 GND.n10 GND.t2 854.365
R15 GND.n10 GND.n0 796.268
R16 GND.n8 GND.n6 792.851
R17 GND.n6 GND.n4 615.143
R18 GND.n2 GND.n0 615.143
R19 GND.n4 GND.t0 239.222
R20 GND.n2 GND.t4 239.222
R21 GND.n13 GND.n12 5.07264
R22 GND.n5 GND.n1 5.05818
R23 GND.n7 GND.n1 4.5005
R24 GND.n12 GND.n11 4.5005
R25 GND.n5 GND.t1 2.17407
R26 GND.n7 GND.t7 2.17389
R27 GND.n11 GND.t3 2.17333
R28 GND.n13 GND.t5 2.17314
R29 GND.n11 GND.n10 2.09407
R30 GND.n8 GND.n7 2.09352
R31 GND.n6 GND.n5 2.09333
R32 GND GND.n0 2.09277
R33 GND.n12 GND.n1 1.97889
R34 GND GND.n13 0.0019876
R35 Q.n2 Q.t4 56.0619
R36 Q.n1 Q.t3 55.9719
R37 Q.n2 Q.t0 4.38208
R38 Q.n1 Q.n0 3.62303
R39 Q.n0 Q.t2 3.0907
R40 Q.n0 Q.t1 2.0905
R41 Q Q.n1 0.108263
R42 Q Q.n2 0.0407632
R43 S S.t0 55.9802
R44 R R.t0 55.985
R45 VDD.n0 VDD.t2 311.146
R46 VDD.n1 VDD.t0 311.132
R47 VDD.n1 VDD.n0 11.0135
R48 VDD.n0 VDD.t3 2.10463
R49 VDD.n1 VDD.t1 2.0905
R50 VDD VDD.n1 0.058473
C0 Qn Q 1.62575f
C1 Q R 0.037842f
C2 Qn S 0.043472f
C3 VDD Q 1.16543f
C4 Qn VDD 0.395392f
C5 R GND 0.256344f
C6 S GND 0.255548f
C7 Q GND 1.65547f
C8 Qn GND 2.41023f
C9 VDD GND 4.11473f
.ends

