* NGSPICE file created from user_proj_sarlogic.ext - technology: gf180mcuD

.subckt user_proj_sarlogic CLK SC SDAC[0] SDAC[1] SDAC[2] SDAC[3] SDAC[4] SDAC[5] SDAC[6] SDAC[7] SDAC[8] XRST COMP_CLK COMP_OUT DIGITAL_OUT vccd1 vssd1
X0 vssd1 a_16569_5984 a_19300_10744 vssd1 nfet_06v0 ad=0.2344p pd=1.56u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1 vccd1 a_24876_3160 a_24976_3608 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2 a_31465_5512 a_29604_9880 vccd1 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X3 a_35424_5644 a_34420_6040 a_35220_5644 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X4 a_13964_7168 a_13656_7212 vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X5 a_6956_11351 a_6868_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X6 a_2588_10216 a_2500_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X7 vccd1 a_11279_7864 a_15492_9521 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X8 a_21852_4076 a_21752_4032 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X9 vccd1 a_24976_3608 SDAC[5] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X10 a_3668_4076 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X11 vssd1 a_15324_6608 a_13496_6366 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X12 a_18268_11784 a_18180_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X13 a_30387_6744 a_27935_4728 a_30199_6744 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X14 a_11279_7864 a_12969_9040 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X15 a_11560_5600 a_2468_4822 a_13572_5176 vccd1 pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X16 a_33096_7124 a_32381_11802 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X17 vccd1 a_16365_5984 a_17456_7080 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X18 a_26564_5176 a_17228_3197 vccd1 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X19 a_23107_5557 a_17640_7564 a_23127_6040 vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X20 a_9385_7952 a_8968_7996 a_9761_7996 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X21 vssd1 a_23756_7080 a_27924_6340 vssd1 nfet_06v0 ad=0.2911p pd=1.53u as=0.3608p ps=2.52u w=0.82u l=0.6u
X22 vccd1 a_5724_10216 a_5636_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X23 vccd1 a_21180_4416 a_25796_9176 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X24 vssd1 CLK a_21392_8392 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X25 vccd1 a_2140_11351 a_2052_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X26 a_17696_4059 a_17284_4472 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X27 a_31341_5557 a_31241_5512 a_30725_5557 vccd1 pfet_06v0 ad=0.37665p pd=1.835u as=0.37665p ps=1.835u w=1.215u l=0.5u
X28 a_16588_11351 a_16500_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X29 a_12992_3988 a_12892_3944 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X30 a_8076_9783 a_7988_9880 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X31 vssd1 a_1908_4118 a_18704_4476 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X32 a_23687_11620 a_23231_11044 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X33 a_30792_9880 a_30240_9880 a_30588_9880 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X34 a_4964_3608 a_4516_3249 vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X35 a_13529_5904 a_13112_6044 a_13905_6044 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X36 vccd1 a_34028_3160 a_32236_3160 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X37 a_11320_6428 a_9520_6744 a_10380_6695 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X38 a_14876_9477 a_18940_7080 a_19089_6744 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X39 a_3528_7612 a_2688_7195 a_3240_7212 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
D0 vssd1 a_2468_3254 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X40 vccd1 a_13900_4728 a_11560_5600 vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X41 a_22560_4292 a_25312_5556 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X42 a_28460_10216 a_28372_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X43 vccd1 a_21392_8392 a_15324_6608 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X44 a_22868_4772 a_21871_5250 vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X45 vssd1 a_35708_9001 SC vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X46 a_19028_5308 a_16108_3228 a_18768_5308 vccd1 pfet_06v0 ad=0.1736p pd=1.18u as=0.224p ps=1.36u w=0.56u l=0.5u
X47 a_24555_7608 a_24435_7098 a_23980_7438 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X48 vccd1 a_17228_3197 a_21871_6818 vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X49 a_3260_8780 a_3140_3272 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X50 vccd1 a_22560_4292 a_35737_4428 vccd1 pfet_06v0 ad=0.4149p pd=2.65u as=0.1521p ps=1.105u w=0.585u l=0.5u
X51 a_14420_4076 a_13252_4472 a_14216_4076 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X52 a_32977_3989 a_27935_4728 a_29772_4773 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X53 a_7050_7124 a_6426_7124 a_6882_7124 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X54 SDAC[0] a_9408_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X55 a_4905_7472 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X56 a_13116_11784 a_13028_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X57 a_27029_10030 a_26909_9432 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X58 a_7924_8312 a_6756_7991 a_7720_8312 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X59 a_7315_3160 a_7645_3160 a_7765_3204 vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X60 a_17416_6016 a_17676_5512 vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
D1 vssd1 a_1908_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X61 vssd1 a_15324_6608 a_27776_7124 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X62 a_32481_11846 a_32381_11802 vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X63 a_35916_7168 a_35608_7212 vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X64 a_22289_6340 a_17004_3197 a_22085_6340 vssd1 nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X65 a_18836_7642 a_16365_5984 vssd1 vssd1 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X66 a_11003_7699 a_10527_7124 a_10751_7146 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X67 a_11123_4381 a_11453_4453 a_11573_4563 vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X68 a_4905_7472 a_4488_7612 a_5281_7612 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X69 vccd1 a_23868_11784 a_23780_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X70 a_22636_11351 a_22548_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X71 a_23751_10030 a_23295_10052 a_23519_9476 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X72 a_11436_11351 a_11348_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X73 vssd1 a_27935_4728 a_33593_4472 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X74 vssd1 a_18403_5949 a_14975_4728 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X75 a_22000_9432 a_19361_6296 vccd1 vccd1 pfet_06v0 ad=0.2486p pd=2.01u as=0.35315p ps=1.96u w=0.565u l=0.5u
X76 a_5713_6744 a_5797_6296 a_5733_6340 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X77 a_19432_8692 a_18828_9199 a_19432_9176 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X78 vccd1 a_16364_6296 a_14567_4728 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X79 a_37904_7864 a_26723_10216 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.2344p ps=1.56u w=0.36u l=0.6u
X80 a_30913_5557 a_20609_5176 a_30725_5557 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X81 a_11304_8780 a_10340_9176 a_11100_8780 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
D2 a_3364_4822 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X82 vccd1 a_12579_10653 a_11740_9500 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X83 vssd1 a_21180_4416 a_34644_7608 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X84 a_3932_11784 a_3844_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X85 vccd1 a_12172_5600 a_12068_5644 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X86 vccd1 a_30723_9085 a_28527_4728 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X87 a_35708_9001 a_37500_9006 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X88 vssd1 a_20096_10688 a_18940_7080 vssd1 nfet_06v0 ad=0.2344p pd=1.56u as=0.3608p ps=2.52u w=0.82u l=0.6u
X89 a_10276_6744 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X90 a_23932_6695 a_23624_6744 vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X91 a_13664_4059 a_13252_4472 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X92 a_14470_7908 a_13994_8484 a_14198_8402 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
D3 vssd1 a_2916_4822 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X93 vccd1 a_28428_3160 SDAC[6] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X94 a_19040_7124 a_18940_7080 a_18836_7124 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X95 vccd1 a_25312_5556 a_22560_4292 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X96 a_15324_6608 a_21392_8392 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X97 a_3772_4032 a_3464_4076 vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X98 a_13564_11784 a_13476_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X99 vssd1 a_15553_5512 a_17640_7564 vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.1248p ps=1u w=0.48u l=0.6u
X100 a_2356_4118 a_13496_6366 vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X101 vssd1 a_18536_10720 a_15383_8679 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X102 vccd1 a_17820_10216 a_17732_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X103 vssd1 a_28540_9500 a_26456_8736 vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X104 vccd1 a_31561_4336 a_31456_4476 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
D4 vssd1 XRST diode_nd2ps_06v0 pj=1.86u area=0.2052p
X105 a_18403_5949 a_18733_6021 a_18853_5578 vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X106 vccd1 a_11123_4381 a_8479_5996 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X107 vccd1 a_1772_7864 DIGITAL_OUT vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X108 a_15464_4476 a_13664_4059 a_14524_4032 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X109 a_17864_8648 a_17456_8648 a_18244_8692 vccd1 pfet_06v0 ad=0.2464p pd=2u as=0.1456p ps=1.08u w=0.56u l=0.5u
X110 vccd1 a_26241_7564 a_23756_7080 vccd1 pfet_06v0 ad=0.38705p pd=2.08u as=0.5368p ps=3.32u w=1.22u l=0.5u
X111 vssd1 a_26241_7564 a_23756_7080 vssd1 nfet_06v0 ad=0.2288p pd=1.58u as=0.3608p ps=2.52u w=0.82u l=0.6u
X112 vccd1 a_32236_3160 SDAC[7] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X113 a_2140_6647 a_2052_6744 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X114 a_13104_7195 a_12692_7608 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X115 a_14216_4076 a_13252_4472 a_14012_4076 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X116 a_11884_11351 a_11796_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X117 vssd1 a_31561_4336 a_31456_4476 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X118 vssd1 a_12580_3608 a_15568_5176 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X119 vssd1 a_36972_7864 a_36044_12281 vssd1 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X120 a_32680_6799 a_32384_6384 a_31623_6564 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.25375p ps=1.51u w=0.505u l=0.5u
X121 a_9644_11351 a_9556_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X122 vccd1 a_35708_9001 SC vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X123 a_13900_11351 a_13812_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X124 a_5276_10216 a_5188_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D5 a_1908_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X125 vccd1 a_21852_10216 a_21764_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X126 vssd1 CLK a_21392_8392 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X127 vccd1 a_18354_6296 a_18474_6916 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X128 vssd1 a_2356_4118 a_7652_4855 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X129 a_23932_6695 a_23624_6744 vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X130 a_19052_8648 a_19300_10744 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2344p ps=1.56u w=0.82u l=0.6u
X131 a_8968_7996 a_6756_7991 a_8028_8263 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X132 vccd1 a_8412_10216 a_8324_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X133 a_37168_10748 a_34644_10744 a_36856_10748 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X134 vccd1 a_21392_8392 a_15324_6608 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X135 a_13533_10792 a_10787_8312 vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X136 a_30723_9085 a_31053_9157 a_31173_9267 vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
D6 vssd1 a_3364_4822 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X137 a_37513_4416 a_36609_4476 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.14985p ps=1.145u w=0.405u l=0.6u
X138 vssd1 a_16108_3228 a_6252_7864 vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.1248p ps=1u w=0.48u l=0.6u
X139 a_21203_7517 a_21533_7589 a_21653_7699 vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
D7 vssd1 a_2356_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X140 SDAC[0] a_9408_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X141 a_28463_4773 a_2916_4822 a_27452_4796 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X142 vccd1 a_2916_4822 a_10599_8312 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X143 vssd1 a_9385_7952 a_9280_7996 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X144 a_4480_6044 a_4332_5600 a_4312_6044 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X145 a_32501_12312 a_32381_11802 vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X146 vccd1 a_1692_9783 a_1604_9880 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X147 a_36680_3205 a_30981_5996 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X148 SDAC[2] a_15568_5176 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X149 vccd1 a_1692_6647 a_1604_6744 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X150 vssd1 a_22000_9432 a_21404_3160 vssd1 nfet_06v0 ad=0.2344p pd=1.56u as=0.3608p ps=2.52u w=0.82u l=0.6u
X151 vccd1 a_1692_3511 a_1604_3608 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X152 a_27753_4336 a_22560_4292 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X153 a_27671_10282 a_27215_10260 a_27439_10282 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X154 vccd1 a_6252_7864 a_15483_8723 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X155 SDAC[5] a_24976_3608 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X156 a_32236_3160 a_34028_3160 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X157 a_29739_6744 a_29075_6875 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2288p ps=1.58u w=0.82u l=0.6u
X158 a_37513_4416 a_36609_4476 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.3276p ps=1.62u w=0.78u l=0.5u
X159 a_21180_4416 a_27776_7124 vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X160 SDAC[2] a_15568_5176 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X161 a_30163_7864 a_30493_7864 a_30613_7908 vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X162 a_18793_9520 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X163 a_21871_6818 a_17640_7564 a_22289_6340 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
X164 vccd1 a_15356_11784 a_15268_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D8 vssd1 CLK diode_nd2ps_06v0 pj=1.86u area=0.2052p
X165 vccd1 a_21180_4416 a_34420_4472 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X166 a_9408_3608 a_7884_8692 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X167 a_7203_6296 a_7533_6296 a_7653_6340 vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
D9 vssd1 a_2468_3254 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X168 SC a_35708_9001 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X169 vccd1 a_22560_4292 a_35737_5996 vccd1 pfet_06v0 ad=0.4149p pd=2.65u as=0.1521p ps=1.105u w=0.585u l=0.5u
X170 vccd1 a_8860_10216 a_8772_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D10 vssd1 a_2468_3254 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X171 a_21392_8392 CLK vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X172 a_26356_10260 a_25908_10791 vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X173 vccd1 a_2468_3254 a_6372_8312 vccd1 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X174 a_28084_5644 a_22560_4292 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X175 a_25368_10720 a_20868_5556 vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X176 a_35210_9476 a_35090_9432 vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X177 vssd1 a_18828_9199 a_19656_9176 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X178 a_23828_6744 a_22660_6423 a_23624_6744 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X179 a_36609_4476 a_34420_4472 a_35737_4428 vccd1 pfet_06v0 ad=0.1079p pd=0.935u as=0.27805p ps=2.17u w=0.415u l=0.5u
X180 a_18388_4728 a_17640_7564 vssd1 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.104p ps=0.92u w=0.4u l=0.6u
X181 a_24097_4476 a_22560_4292 vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X182 vccd1 a_2356_4118 a_16164_9559 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X183 a_4024_5644 a_3472_5627 a_3820_5644 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X184 a_10871_7864 a_10751_7146 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X185 a_35708_9001 a_37500_9006 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X186 vssd1 a_30723_9085 a_28527_4728 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X187 a_14533_5557 a_13529_5904 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X188 a_4760_6341 a_5020_6341 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X189 a_20289_4476 a_1908_4118 vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X190 vssd1 a_1908_4118 a_17584_9564 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X191 COMP_CLK a_33916_11000 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X192 vssd1 a_19656_7909 a_17004_3197 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X193 vssd1 a_35708_11000 a_33916_11000 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X194 vccd1 a_1692_10216 a_1604_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X195 a_3619_4728 a_3949_4728 a_4069_5326 vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X196 vccd1 a_33461_9477 a_37780_9568 vccd1 pfet_06v0 ad=0.35315p pd=1.96u as=0.2486p ps=2.01u w=0.565u l=0.5u
X197 a_23304_4476 a_21092_4472 a_22364_4032 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X198 a_16252_11784 a_16164_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X199 a_27358_11850 a_26902_12404 a_27126_11850 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X200 vccd1 a_37912_4773 a_37196_11045 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X201 a_7884_8692 a_7428_9176 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.35315p ps=1.96u w=1.22u l=0.5u
X202 a_18704_4476 a_18556_4032 a_18536_4476 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X203 a_20096_10688 a_19916_7909 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.2344p ps=1.56u w=0.36u l=0.6u
X204 vssd1 a_17456_8648 a_17864_8648 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X205 vccd1 a_25100_11351 a_25012_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X206 vccd1 a_10204_11784 a_10116_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X207 vssd1 a_26579_9432 a_24435_7098 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X208 vccd1 a_1692_8648 a_1604_8692 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X209 a_36833_4476 a_34420_4472 a_36609_4476 vssd1 nfet_06v0 ad=0.2898p pd=2.33u as=93.59999f ps=0.88u w=0.36u l=0.6u
X210 vccd1 a_1692_5512 a_1604_5556 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X211 a_4800_7612 a_2276_7608 a_4488_7612 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X212 a_14533_5557 a_13529_5904 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X213 a_32995_11784 a_37273_10608 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X214 vccd1 a_15030_7908 a_15486_8462 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X215 a_23721_4336 a_22560_4292 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X216 a_20411_6760 a_17004_3197 a_20615_6340 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X217 a_5505_9180 a_1908_4118 vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X218 vccd1 a_5612_9783 a_5524_9880 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X219 vssd1 a_15568_5176 SDAC[2] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X220 a_11285_4773 a_10281_4816 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X221 a_18828_9199 a_20403_7098 vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X222 a_31117_7864 a_31509_7864 vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X223 a_25866_11828 a_25242_11828 a_25718_12404 vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X224 a_34412_9176 a_34292_8648 a_34144_9238 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.2569p ps=1.56u w=0.82u l=0.6u
X225 a_31117_4728 a_23599_5996 vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X226 a_6882_7124 a_6426_7124 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X227 a_15568_5176 a_12580_3608 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X228 vccd1 a_17820_11784 a_17732_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X229 a_7765_3204 a_7645_3160 vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X230 a_4228_5644 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X231 a_23420_6744 a_23320_6574 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X232 vccd1 a_24540_10216 a_24452_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X233 a_4712_4476 a_2500_4472 a_3772_4032 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X234 vssd1 a_1908_4118 a_12320_6044 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X235 vssd1 a_35708_9001 SC vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X236 a_11573_4563 a_11453_4453 vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X237 vssd1 a_33094_5892 a_2468_3254 vssd1 nfet_06v0 ad=0.2911p pd=1.53u as=0.2132p ps=1.34u w=0.82u l=0.6u
X238 vccd1 a_34888_9152 a_32404_7864 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X239 a_23616_4476 a_21504_4059 a_23304_4476 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X240 a_24675_4728 a_25005_4728 a_25125_5326 vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X241 vssd1 a_32457_9520 a_32352_9564 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X242 a_11100_11784 a_11012_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X243 a_18648_4748 a_16365_5984 vssd1 vssd1 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X244 a_16512_9120 a_16325_7125 vccd1 vccd1 pfet_06v0 ad=0.2486p pd=2.01u as=0.35315p ps=1.96u w=0.565u l=0.5u
X245 a_3696_3608 a_3596_3228 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X246 vccd1 a_9408_3608 SDAC[0] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X247 SDAC[0] a_9408_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X248 a_16824_9710 a_17456_8648 a_17368_8692 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X249 vssd1 a_2468_3254 a_24555_7608 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X250 a_11760_9180 a_11612_8736 a_11592_9180 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X251 a_11312_5627 a_10900_6040 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X252 a_7168_8312 a_6756_7991 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X253 vccd1 a_32872_6686 a_32680_6799 vccd1 pfet_06v0 ad=0.2222p pd=1.89u as=0.2424p ps=1.465u w=0.505u l=0.5u
X254 vssd1 a_27924_6340 a_2468_4822 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X255 a_27935_4728 a_28040_7944 a_30778_7124 vccd1 pfet_06v0 ad=0.3477p pd=1.79u as=0.4087p ps=1.89u w=1.22u l=0.5u
X256 vccd1 a_6396_11784 a_6308_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X257 vccd1 a_2356_4118 a_2500_9176 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X258 a_33916_11000 a_35708_11000 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X259 vssd1 a_32236_3160 SDAC[7] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X260 vccd1 a_10652_11784 a_10564_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X261 a_30240_9880 a_29828_9559 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X262 a_35220_5644 a_35100_5996 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X263 vssd1 a_11737_6384 a_11632_6428 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X264 a_33461_9477 a_32457_9520 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X265 a_35677_4076 a_34420_4472 a_35424_4076 vccd1 pfet_06v0 ad=0.101p pd=0.905u as=0.19315p ps=1.27u w=0.505u l=0.5u
X266 a_10983_7146 a_10527_7124 a_10751_7146 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X267 vccd1 a_31750_7460 a_2916_4822 vccd1 pfet_06v0 ad=0.4941p pd=2.03u as=0.3782p ps=1.84u w=1.22u l=0.5u
X268 vssd1 a_31750_7460 a_2916_4822 vssd1 nfet_06v0 ad=0.2911p pd=1.53u as=0.2132p ps=1.34u w=0.82u l=0.6u
D11 vssd1 a_3364_4822 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X269 vssd1 a_32381_11802 a_33992_7608 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X270 vccd1 XRST a_4516_3249 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X271 a_12892_3944 a_3364_4822 a_14295_5176 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
D12 a_2356_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X272 vccd1 a_32384_6384 a_32279_6755 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X273 a_13496_6366 a_15324_6608 vssd1 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X274 a_33768_7124 a_32381_11802 a_33768_7608 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3172p ps=1.74u w=1.22u l=0.5u
X275 vssd1 a_1908_4118 a_3696_7612 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X276 vccd1 a_2356_4118 a_2276_7608 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X277 vccd1 a_3036_9783 a_2948_9880 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X278 a_32236_3160 a_34028_3160 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X279 a_19447_5176 a_20127_4728 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X280 vccd1 a_6496_3988 a_1908_4118 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X281 a_24872_6428 a_22660_6423 a_23932_6695 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X282 a_27753_4336 a_27336_4476 a_28129_4476 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X283 a_21180_4416 a_27776_7124 vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X284 a_31453_10792 a_29244_9477 vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X285 a_25884_4076 a_25784_4032 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X286 a_36081_6044 a_35424_5644 vssd1 vssd1 nfet_06v0 ad=86.399994f pd=0.84u as=93.59999f ps=0.88u w=0.36u l=0.6u
X287 a_33339_12404 a_32863_11828 vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X288 a_9408_3608 a_7884_8692 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X289 a_5020_6341 a_6133_3989 a_6887_4773 vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X290 vssd1 a_2356_4118 a_17284_4472 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X291 a_18853_5578 a_18733_6021 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X292 a_15321_7472 a_14904_7612 a_15697_7612 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X293 a_20844_8780 a_19432_9176 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X294 a_24115_5557 a_20868_5556 a_23927_5557 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X295 a_27776_7124 a_15324_6608 vssd1 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X296 a_7292_11784 a_7204_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X297 a_36008_3205 a_35428_3608 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X298 a_18388_4728 a_18648_4748 vssd1 vssd1 nfet_06v0 ad=0.14p pd=1.1u as=0.224p ps=1.52u w=0.4u l=0.6u
X299 a_4257_6744 a_4341_6296 a_4277_6340 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X300 a_23652_7608 a_23756_7080 a_23652_7124 vccd1 pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X301 a_15324_6608 a_21392_8392 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X302 SDAC[1] a_13216_3608 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X303 a_15940_9880 a_15492_9521 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X304 SC a_35708_9001 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X305 a_13900_4728 a_14567_4728 vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X306 a_3696_3608 a_3596_3228 vssd1 vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X307 vssd1 a_37513_4416 a_37465_4472 vssd1 nfet_06v0 ad=0.14985p pd=1.145u as=48.6f ps=0.645u w=0.405u l=0.6u
X308 a_26487_11620 a_26031_11044 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X309 vssd1 a_21203_5949 a_20127_4728 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X310 vssd1 a_9408_3608 SDAC[0] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X311 a_19357_6088 a_12220_3205 vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
D13 vssd1 a_1908_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X312 a_2588_11351 a_2500_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X313 a_12579_10653 a_12909_10725 a_13029_10282 vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X314 a_18474_6916 a_18354_6296 a_17730_6296 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X315 a_37273_7472 a_36856_7612 a_37649_7612 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X316 vccd1 a_32236_3160 SDAC[7] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X317 vssd1 a_17456_8648 a_20523_7608 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X318 a_11660_5644 a_11560_5600 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X319 a_30163_7864 a_30493_7864 a_30613_8462 vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X320 vccd1 a_29356_10216 a_29268_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X321 vccd1 a_22076_11784 a_21988_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X322 a_30163_4728 a_30493_4728 a_30613_5326 vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X323 vccd1 a_11740_9500 a_11000_8736 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X324 vccd1 a_15568_5176 SDAC[2] vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X325 a_37273_7472 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X326 a_9084_9783 a_8996_9880 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X327 vccd1 a_32507_4728 a_30981_5996 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X328 vccd1 a_4380_10216 a_4292_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X329 a_5972_3608 a_5524_3249 vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
D14 a_2356_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X330 a_35737_5996 a_22560_4292 a_36081_6044 vssd1 nfet_06v0 ad=0.1989p pd=1.465u as=86.399994f ps=0.84u w=0.36u l=0.6u
X331 vccd1 a_6508_11351 a_6420_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X332 a_37273_10608 a_22560_4292 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X333 a_31173_9267 a_31053_9157 vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X334 vccd1 a_6133_8693 a_6140_4728 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X335 vccd1 a_15464_4476 a_15881_4336 vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X336 a_33766_10596 a_33461_9477 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2911p ps=1.53u w=0.82u l=0.6u
X337 a_27236_6340 a_23756_7080 a_27236_6744 vccd1 pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X338 a_22344_4476 a_21504_4059 a_22056_4076 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X339 a_21653_7699 a_21533_7589 vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X340 vccd1 a_24976_3608 SDAC[5] vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X341 a_32457_9520 a_22560_4292 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X342 vccd1 a_27564_6296 a_27236_6340 vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X343 a_34104_6384 a_30387_6744 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X344 a_5797_6296 a_8310_7146 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X345 a_2140_11784 a_2052_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X346 vssd1 a_15568_5176 SDAC[2] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X347 vssd1 a_27215_10260 a_27691_10835 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X348 a_11100_8780 a_11000_8736 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X349 a_4312_6044 a_3472_5627 a_4024_5644 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X350 a_11508_8780 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X351 a_30913_5557 a_31465_5512 vssd1 vssd1 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X352 a_24092_10216 a_24004_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X353 a_24249_9880 a_23519_9476 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X354 vccd1 a_37500_9006 a_35708_9001 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X355 a_3036_7212 a_2936_7168 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X356 vssd1 a_14616_9477 a_12188_7864 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X357 a_21203_5949 a_21533_6021 a_21653_5578 vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X358 vccd1 a_1692_11784 a_1604_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X359 DIGITAL_OUT a_1772_7864 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X360 a_4828_10216 a_4740_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X361 vssd1 a_32380_5870 a_31844_6040 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X362 a_16485_6040 a_16365_5984 a_16291_6040 vssd1 nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X363 a_31148_11784 a_31060_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D15 vssd1 a_2356_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X364 a_9385_7952 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
D16 vssd1 a_2916_4822 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X365 vssd1 a_33766_10596 a_28040_7944 vssd1 nfet_06v0 ad=0.2911p pd=1.53u as=0.2132p ps=1.34u w=0.82u l=0.6u
X366 vccd1 a_21392_8392 a_15324_6608 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X367 a_36084_6377 a_28428_7944 a_36064_6744 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X368 a_37273_10608 a_36856_10748 a_37649_10748 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X369 vccd1 a_9408_3608 SDAC[0] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X370 a_29176_7909 a_26513_7471 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X371 a_30613_7908 a_30493_7864 vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X372 vssd1 a_28527_4728 a_28463_4773 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X373 vccd1 a_32457_9520 a_32352_9564 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X374 a_9632_5556 a_9532_5512 vssd1 vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X375 a_7653_6340 a_7533_6296 vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X376 a_31456_4476 a_28932_4472 a_31144_4476 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X377 a_21292_11351 a_21204_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X378 a_12556_4773 a_15553_5512 a_15057_5557 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X379 a_10092_11351 a_10004_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X380 vssd1 a_31304_3205 a_30220_3160 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X381 vssd1 a_17864_7080 a_13352_7168 vssd1 nfet_06v0 ad=0.218p pd=1.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X382 SDAC[7] a_32236_3160 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X383 a_19357_6088 a_12220_3205 vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X384 vccd1 a_6956_11351 a_6868_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X385 vssd1 a_12244_5176 a_13216_3608 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X386 a_17676_5512 a_3364_4822 a_19447_5176 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X387 vccd1 a_24540_11784 a_24452_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X388 vccd1 a_30204_4032 a_30100_4076 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X389 vccd1 a_3484_9783 a_3396_9880 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X390 a_31237_7908 a_31117_7864 a_30493_7864 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X391 a_23855_11620 a_23231_11044 a_23687_11620 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X392 a_5129_4336 a_4712_4476 a_5505_4476 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X393 vccd1 a_28008_9180 a_28425_9040 vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X394 a_19524_11448 a_19076_11089 vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X395 vccd1 a_23756_7080 a_27924_6340 vccd1 pfet_06v0 ad=0.4941p pd=2.03u as=0.5368p ps=3.32u w=1.22u l=0.5u
X396 a_21392_8392 CLK vssd1 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X397 vccd1 a_16588_11351 a_16500_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X398 a_17584_9564 a_17436_9831 a_17416_9564 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X399 a_34104_5118 a_33616_4816 a_34364_5176 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X400 vccd1 a_15321_7472 a_15216_7612 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X401 a_11003_9476 a_10871_7864 a_10428_5870 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X402 vccd1 a_15568_5176 SDAC[2] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X403 a_10527_7124 a_9903_7124 a_10379_7700 vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X404 a_27900_11351 a_27812_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X405 a_36884_9880 a_33461_9477 a_36268_12281 vccd1 pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X406 a_23363_11000 a_37513_4416 vccd1 vccd1 pfet_06v0 ad=0.6561p pd=3.51u as=0.5346p ps=3.31u w=1.215u l=0.5u
X407 vccd1 a_17318_6562 a_17418_6916 vccd1 pfet_06v0 ad=0.1656p pd=1.28u as=61.199993f ps=0.7u w=0.36u l=0.5u
X408 a_35428_3608 a_34980_3249 vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X409 vccd1 a_14908_11784 a_14820_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X410 vssd1 a_25368_10720 a_15737_5996 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X411 vssd1 a_21180_4416 a_34644_10744 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X412 a_4712_9180 a_2912_8763 a_3772_8736 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X413 vccd1 a_10428_10216 a_10340_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X414 vssd1 a_15321_7472 a_15216_7612 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X415 a_22713_9040 a_22296_9180 a_23089_9180 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X416 a_15486_8462 a_15030_7908 a_15254_7908 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X417 a_6036_4772 a_2468_4822 a_4965_4728 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
D17 a_2916_4822 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X418 a_32481_11846 a_32565_12256 a_32501_12312 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X419 vssd1 a_9408_3608 SDAC[0] vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X420 SDAC[0] a_9408_3608 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X421 a_27847_5176 a_28119_4728 a_27452_4796 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X422 a_33284_7124 a_32381_11802 a_33096_7124 vccd1 pfet_06v0 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.5u
X423 a_25289_6384 a_24872_6428 a_25665_6428 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X424 vccd1 a_37273_7472 a_37168_7612 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X425 a_12580_3608 a_12132_3249 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X426 vssd1 a_18940_7080 a_18836_7642 vssd1 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X427 vccd1 a_22636_11351 a_22548_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X428 a_34832_5627 a_34420_6040 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X429 a_33500_9006 a_32404_7864 a_34069_6040 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X430 vssd1 a_37273_7472 a_37168_7612 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X431 vccd1 a_11436_11351 a_11348_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X432 vssd1 a_12580_3608 a_15568_5176 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
D18 vssd1 a_2356_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X433 a_20868_5556 a_20420_6087 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X434 a_15804_11784 a_15716_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X435 vccd1 a_35708_9001 SC vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X436 vssd1 a_17318_6562 a_17458_6340 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X437 a_11592_9180 a_10752_8763 a_11304_8780 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X438 vssd1 CLK a_21392_8392 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X439 a_29263_6875 a_26456_8736 a_29075_6875 vccd1 pfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.5u
X440 vssd1 a_21203_7517 a_20403_7098 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X441 a_12320_6044 a_12172_5600 a_12152_6044 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X442 vccd1 a_21203_7517 a_20403_7098 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X443 vccd1 a_26396_4032 a_26292_4076 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X444 vccd1 a_10281_4816 a_10176_4860 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X445 a_35100_5996 a_32481_11846 a_36884_6340 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X446 vssd1 a_31465_5512 a_34412_9176 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X447 a_28757_3989 a_27753_4336 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X448 a_17332_9880 a_16164_9559 a_17128_9880 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X449 a_3472_5627 a_3060_6040 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X450 SDAC[8] a_33916_7864 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X451 vccd1 a_10876_10216 a_10788_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X452 a_3696_7612 a_3548_7168 a_3528_7612 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X453 a_36609_4476 a_34832_4059 a_35737_4428 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1989p ps=1.465u w=0.36u l=0.6u
X454 vccd1 a_19768_7584 a_18236_7864 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X455 vccd1 a_4380_11784 a_4292_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X456 vccd1 a_21356_8736 a_21252_8780 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X457 vccd1 a_13964_7168 a_13860_7212 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X458 vccd1 a_21392_8392 a_15324_6608 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X459 a_7516_10216 a_7428_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X460 vssd1 a_37500_9006 a_35708_9001 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X461 vssd1 a_33916_11000 COMP_CLK vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X462 a_1908_4118 a_6496_3988 vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X463 a_26241_7564 a_2468_3254 a_26633_7124 vccd1 pfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.5u
X464 vccd1 a_37912_11045 a_35708_11000 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X465 a_30407_6341 a_27935_4728 vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X466 a_28757_3989 a_27753_4336 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X467 a_36044_12281 a_36972_7864 a_37968_6744 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X468 vssd1 a_37912_12288 a_16108_3228 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X469 a_7416_8142 a_9980_5870 a_9892_6040 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X470 a_22085_6340 a_17228_3197 a_21891_6340 vssd1 nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
D19 vssd1 a_1908_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
D20 a_2356_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X471 a_35812_10348 a_22560_4292 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X472 vccd1 a_2140_9783 a_2052_9880 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D21 a_2356_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X473 a_17864_8648 a_16365_5984 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.218p ps=1.52u w=0.36u l=0.6u
X474 a_8412_5176 a_3696_3608 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X475 vccd1 a_2140_6647 a_2052_6744 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X476 a_35608_10348 a_34644_10744 a_35404_10348 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X477 vccd1 a_28425_9040 a_28320_9180 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X478 vccd1 a_11884_11351 a_11796_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X479 vccd1 a_5948_11784 a_5860_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X480 vccd1 a_9644_11351 a_9556_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X481 a_19916_7909 a_22713_9040 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X482 vccd1 a_29128_6044 a_29545_5904 vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X483 a_19705_6341 a_18940_7080 a_14876_9477 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X484 a_33916_11000 a_35708_11000 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X485 SDAC[6] a_28428_3160 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X486 a_15940_9880 a_15492_9521 vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X487 vccd1 a_5129_4336 a_5024_4476 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X488 vccd1 a_13900_11351 a_13812_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X489 a_37465_4472 a_22560_4292 a_36833_4476 vssd1 nfet_06v0 ad=48.6f pd=0.645u as=0.3123p ps=2.38u w=0.405u l=0.6u
X490 a_4760_6341 a_5020_6341 vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X491 vccd1 a_31117_7864 a_31237_8484 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X492 a_37912_12288 COMP_OUT vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X493 vccd1 a_31117_4728 a_31237_5348 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X494 a_17456_7080 a_18940_7080 a_18935_7908 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X495 a_14420_4076 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X496 a_13905_6044 a_1908_4118 vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X497 a_10380_6695 a_10072_6744 vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X498 vccd1 a_1772_7864 DIGITAL_OUT vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X499 a_10072_6744 a_9520_6744 a_9868_6744 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X500 a_25536_4059 a_25124_4472 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X501 a_25548_11351 a_25460_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X502 a_14348_11351 a_14260_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X503 a_7964_10216 a_7876_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X504 vccd1 a_2916_4822 a_6679_5176 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X505 a_8924_5127 a_8616_5176 vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X506 vccd1 a_33916_7864 SDAC[8] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X507 SDAC[0] a_9408_3608 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X508 a_27029_9476 a_26909_9432 vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X509 vccd1 a_20060_11784 a_19972_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X510 vssd1 a_11740_9500 a_11000_8736 vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X511 a_35424_5644 a_34832_5627 a_35220_5644 vccd1 pfet_06v0 ad=0.19315p pd=1.27u as=0.1313p ps=1.025u w=0.505u l=0.5u
X512 a_6844_11784 a_6756_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X513 a_27116_6296 a_26804_7953 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X514 a_2468_4822 a_27924_6340 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2911p ps=1.53u w=0.82u l=0.6u
D22 vssd1 a_2356_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X515 a_13345_9180 a_1908_4118 vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X516 a_36064_6744 a_32381_11802 vccd1 vccd1 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X517 a_2356_4118 a_13496_6366 vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X518 vccd1 a_2356_4118 a_12692_7608 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X519 a_20496_8763 a_20084_9176 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
D23 vssd1 a_2356_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X520 a_22848_5176 a_21871_5250 a_22660_5176 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X521 a_35404_7212 a_27609_11448 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X522 a_31623_6564 a_32384_6384 a_32175_6799 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=94.5f ps=0.885u w=0.36u l=0.6u
X523 vccd1 a_25289_6384 a_25184_6428 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X524 a_25248_9120 a_23599_5996 vccd1 vccd1 pfet_06v0 ad=0.2486p pd=2.01u as=0.35315p ps=1.96u w=0.565u l=0.5u
X525 vssd1 a_1772_7864 DIGITAL_OUT vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X526 a_2916_4822 a_31750_7460 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X527 vccd1 a_19656_7909 a_17004_3197 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X528 a_21653_5578 a_21533_6021 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X529 a_2916_4822 a_31750_7460 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X530 a_13216_3608 a_12244_5176 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X531 a_13496_6366 a_15324_6608 vccd1 vccd1 pfet_06v0 ad=0.2952p pd=1.54u as=0.367p ps=1.92u w=0.82u l=0.5u
X532 vccd1 a_34028_3160 a_32236_3160 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X533 vccd1 a_2140_8648 a_2052_8692 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X534 a_29739_6744 a_29075_6875 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.38705p ps=2.08u w=1.22u l=0.5u
X535 vccd1 a_36268_12281 a_36154_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X536 vccd1 a_35737_4428 a_35677_4076 vccd1 pfet_06v0 ad=0.3975p pd=2.185u as=0.101p ps=0.905u w=0.505u l=0.5u
X537 vccd1 a_31465_5512 a_32380_5870 vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X538 vccd1 a_28908_10216 a_28820_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X539 a_20609_5176 a_6252_7864 a_20629_4772 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X540 a_4573_4728 a_4965_4728 vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X541 a_28160_7988 a_28040_7944 vssd1 vssd1 nfet_06v0 ad=79.799995f pd=0.8u as=0.2424p ps=1.635u w=0.38u l=0.6u
X542 vccd1 a_21628_11784 a_21540_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X543 vccd1 a_21180_4416 a_34644_7608 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X544 a_28428_3160 a_30220_3160 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X545 vssd1 a_7884_8692 a_9408_3608 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X546 a_8157_6296 a_5909_7125 vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X547 vccd1 a_32040_9564 a_32457_9520 vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X548 a_9408_3608 a_7884_8692 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X549 vssd1 a_32872_6686 a_32680_6799 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=0.2007p ps=1.475u w=0.36u l=0.6u
X550 a_13860_7212 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X551 vccd1 a_2356_4118 a_20084_9176 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X552 vccd1 a_3932_10216 a_3844_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X553 DIGITAL_OUT a_1772_7864 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X554 vssd1 a_27935_4728 a_34980_6340 vssd1 nfet_06v0 ad=0.2911p pd=1.53u as=0.3608p ps=2.52u w=0.82u l=0.6u
X555 a_22157_6088 a_19361_6296 vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X556 vccd1 a_3772_4032 a_3668_4076 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X557 a_14796_11351 a_14708_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D24 vssd1 a_2916_4822 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X558 vccd1 a_21180_4416 a_34644_10744 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X559 a_10752_8763 a_10340_9176 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X560 a_17241_7909 a_16325_7125 a_12860_7909 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X561 a_10599_8312 a_10871_7864 a_10787_8312 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
D25 a_16108_3228 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X562 vccd1 a_26902_12404 a_27358_11850 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X563 vssd1 a_22560_4292 a_22512_4476 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X564 a_21504_4059 a_21092_4472 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X565 vccd1 a_4964_3608 a_5524_3249 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X566 a_23644_10216 a_23556_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X567 a_30240_9880 a_29828_9559 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X568 a_22608_9180 a_20084_9176 a_22296_9180 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X569 vccd1 a_31304_3205 a_30220_3160 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X570 a_1908_4118 a_6496_3988 vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X571 a_26293_6341 a_25289_6384 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X572 vccd1 a_24360_9152 a_23200_4728 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X573 SDAC[0] a_9408_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X574 vccd1 a_19357_6088 a_19477_5556 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X575 a_7416_8142 a_2468_4822 a_10100_5556 vccd1 pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X576 a_23624_6744 a_22660_6423 a_23420_6744 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X577 a_22524_11784 a_22436_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X578 vccd1 a_30700_11784 a_30612_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X579 a_17416_9564 a_16576_9880 a_17128_9880 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X580 vccd1 a_4964_3608 a_6496_3988 vccd1 pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X581 vssd1 a_18940_7080 a_18648_4748 vssd1 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X582 a_37912_4773 a_33768_7608 vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X583 vccd1 a_20411_6760 a_22919_5557 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X584 a_13826_8484 a_13370_7908 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X585 a_16325_7125 a_15321_7472 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X586 a_19916_7909 a_22713_9040 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X587 vssd1 a_33616_4816 a_33511_5187 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X588 a_34441_11828 a_33711_11850 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X589 a_10379_7700 a_9903_7124 vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X590 a_37092_7908 a_36972_7864 vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X591 a_26760_8780 a_26208_8763 a_26556_8780 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X592 DIGITAL_OUT a_1772_7864 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
D26 a_2468_3254 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X593 a_22056_4076 a_21092_4472 a_21852_4076 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X594 a_31509_7864 a_2468_4822 a_32052_5556 vccd1 pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X595 a_37912_11045 a_32995_11784 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X596 vssd1 a_1908_4118 a_3920_4476 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X597 a_18452_4076 a_17284_4472 a_18248_4076 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X598 a_5272_6044 a_3472_5627 a_4332_5600 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X599 vccd1 a_29739_6744 a_30199_6744 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X600 SDAC[6] a_28428_3160 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X601 a_29512_4773 a_29772_4773 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X602 SDAC[2] a_15568_5176 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X603 vccd1 a_8636_11784 a_8548_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X604 a_33766_10596 a_33461_9477 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4941p ps=2.03u w=1.22u l=0.5u
X605 a_2356_4118 a_13496_6366 vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.5368p ps=3.32u w=1.22u l=0.5u
X606 a_7404_11351 a_7316_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X607 vssd1 a_23052_7564 a_21752_4032 vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X608 vccd1 a_19496_4476 a_19913_4336 vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X609 vccd1 a_12580_3608 a_15568_5176 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X610 vssd1 a_31241_5512 a_30913_5557 vssd1 nfet_06v0 ad=0.1209p pd=0.985u as=0.21175p ps=1.41u w=0.465u l=0.6u
X611 a_17318_6562 a_17730_6296 a_17850_6340 vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X612 a_26723_10216 a_37273_7472 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X613 vccd1 a_23052_7564 a_21752_4032 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
D27 vssd1 a_2468_3254 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X614 a_35708_9001 a_37500_9006 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X615 a_3036_10216 a_2948_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X616 a_35812_10348 a_34644_10744 a_35608_10348 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X617 a_14503_4773 a_3364_4822 vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X618 vssd1 a_29244_9477 a_29156_9521 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X619 vccd1 a_1772_7864 DIGITAL_OUT vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X620 vccd1 a_32404_7864 a_31465_5512 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X621 vssd1 a_28425_9040 a_28320_9180 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X622 a_2912_4059 a_2500_4472 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X623 a_27776_7124 a_15324_6608 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X624 a_22157_6088 a_19361_6296 vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X625 a_37968_6744 a_32481_11846 vccd1 vccd1 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
D28 a_2916_4822 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X626 a_6440_9152 a_5909_7125 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X627 a_3464_4076 a_2500_4472 a_3260_4076 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X628 a_13104_7195 a_12692_7608 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X629 SDAC[0] a_9408_3608 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X630 vccd1 a_18268_11784 a_18180_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X631 a_26396_4032 a_26088_4076 vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X632 a_17036_11351 a_16948_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X633 vccd1 a_4712_9180 a_5129_9040 vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X634 a_9633_4006 a_2468_3254 vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X635 a_22972_11784 a_22884_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X636 COMP_CLK a_33916_11000 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X637 a_35404_10348 a_35304_10304 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X638 vccd1 a_21180_4416 a_29828_9559 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X639 a_26964_8780 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X640 vccd1 a_27924_6340 a_2468_4822 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X641 a_17458_6340 a_17318_6562 a_16694_6296 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
D29 vssd1 a_2356_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X642 vssd1 a_6496_3988 a_1908_4118 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X643 vccd1 a_12188_7864 a_12084_8312 vccd1 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X644 a_17368_7124 a_17640_7564 a_13352_7168 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X645 a_13352_7168 a_17640_7564 a_17576_7608 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X646 a_21356_8736 a_21048_8780 vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X647 vssd1 a_19357_6088 a_19477_6132 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X648 a_12152_6044 a_11312_5627 a_11864_5644 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
D30 vssd1 a_2468_4822 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X649 a_30588_9880 a_30488_9710 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X650 a_8008_7996 a_7168_8312 a_7720_8312 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X651 a_20431_6340 a_6252_7864 vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
D31 a_2468_3254 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X652 a_28040_7944 a_33766_10596 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X653 a_17696_4059 a_17284_4472 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X654 a_13216_3608 a_12244_5176 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X655 a_13496_6366 a_15324_6608 vccd1 vccd1 pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
D32 vssd1 a_3364_4822 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X656 a_33724_9432 a_34054_9432 a_34174_9476 vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X657 a_13964_7168 a_13656_7212 vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X658 vccd1 a_29545_5904 a_29440_6044 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X659 vssd1 a_18388_4728 a_15329_5996 vssd1 nfet_06v0 ad=0.224p pd=1.52u as=0.3608p ps=2.52u w=0.82u l=0.6u
X660 a_7852_11351 a_7764_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X661 a_37172_4772 a_37500_4728 a_37152_5194 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X662 a_4828_11351 a_4740_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X663 a_9408_3608 a_7884_8692 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X664 vssd1 a_7884_8692 a_9408_3608 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X665 a_14216_4076 a_13664_4059 a_14012_4076 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X666 a_3484_10216 a_3396_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X667 a_25159_7125 a_25839_7564 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X668 a_18836_7642 a_15553_5512 a_19040_7124 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X669 a_19164_11784 a_19076_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X670 vssd1 a_28428_3160 SDAC[6] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X671 a_33616_4816 a_21180_4416 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X672 a_35916_7168 a_35608_7212 vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X673 vccd1 a_29604_9880 a_31465_5512 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X674 a_19496_4476 a_17696_4059 a_18556_4032 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X675 vssd1 a_32507_4728 a_30981_5996 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X676 a_17870_6916 a_17730_6296 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1656p ps=1.28u w=0.36u l=0.5u
X677 a_19169_9564 a_1908_4118 vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X678 a_36972_7864 a_37780_9568 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.35315p ps=1.96u w=1.22u l=0.5u
X679 vccd1 a_13116_11784 a_13028_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X680 vccd1 a_13994_8484 a_14430_8484 vccd1 pfet_06v0 ad=0.1656p pd=1.28u as=61.199993f ps=0.7u w=0.36u l=0.5u
X681 a_26655_11620 a_26031_11044 a_26487_11620 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X682 SDAC[2] a_15568_5176 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
D33 vssd1 a_3364_4822 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X683 a_18248_4076 a_17284_4472 a_18044_4076 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X684 vccd1 a_6620_10216 a_6532_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X685 DIGITAL_OUT a_1772_7864 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X686 vssd1 a_2356_4118 a_12692_7608 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
D34 vssd1 a_1908_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X687 a_17484_11351 a_17396_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X688 vccd1 a_7315_3160 a_4229_3160 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X689 a_4965_4728 a_6140_4728 a_6036_4772 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X690 vssd1 a_4760_6341 a_3228_3228 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X691 a_21180_4416 a_27776_7124 vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X692 a_19432_9176 a_19052_8648 a_19432_8692 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X693 a_31937_4476 a_22560_4292 vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X694 vccd1 a_9408_3608 SDAC[0] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X695 a_13112_6044 a_11312_5627 a_12172_5600 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X696 a_33916_7864 a_35708_7864 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X697 vssd1 a_8269_3160 a_8389_3204 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X698 vccd1 a_2588_11351 a_2500_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X699 a_31237_8484 a_31117_7864 a_30493_7864 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X700 SC a_35708_9001 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X701 a_31237_5348 a_31117_4728 a_30493_4728 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X702 a_37168_7612 a_34644_7608 a_36856_7612 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X703 a_33768_7608 a_32565_12256 a_33768_7124 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X704 a_36856_10748 a_35056_10331 a_35916_10304 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
D35 a_2356_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X705 a_21392_8392 CLK vssd1 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X706 vccd1 a_3932_11784 a_3844_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X707 a_37500_4728 a_37108_11089 vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X708 a_32175_6799 a_31275_6296 vccd1 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.29465p ps=1.74u w=0.505u l=0.5u
X709 vssd1 a_32236_3160 SDAC[7] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X710 a_10281_4816 a_9864_4860 a_10657_4860 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X711 a_28169_10260 a_27439_10282 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X712 a_20844_8780 a_19432_9176 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X713 a_26544_4476 a_26396_4032 a_26376_4476 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X714 vssd1 a_10527_7124 a_11003_7699 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X715 a_14012_11784 a_13924_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X716 a_18751_7908 a_17456_8648 vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X717 SDAC[8] a_33916_7864 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
D36 vssd1 a_1908_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X718 a_6252_7864 a_16108_3228 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X719 vssd1 a_13216_3608 SDAC[1] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X720 a_31304_3205 a_24607_5996 vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X721 a_12579_10653 a_12909_10725 a_13029_10835 vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X722 vccd1 a_30981_5996 a_32977_3989 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X723 a_25159_7125 a_24435_7098 a_23052_7564 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X724 a_26356_10260 a_25908_10791 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X725 a_12552_9180 a_10752_8763 a_11612_8736 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X726 a_18836_7124 a_16365_5984 vccd1 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X727 vssd1 a_16365_5984 a_19705_6341 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X728 vccd1 a_13564_11784 a_13476_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X729 a_12332_11351 a_12244_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X730 vssd1 XRST a_4516_3249 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X731 a_17228_3197 a_20495_6296 vssd1 vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X732 a_19655_4773 a_3364_4822 vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X733 a_27068_8736 a_26760_8780 vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X734 a_25184_6428 a_22660_6423 a_24872_6428 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X735 a_29804_11784 a_29716_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X736 a_32748_7908 a_32404_7864 a_31465_5512 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X737 vccd1 a_15568_5176 SDAC[2] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X738 vccd1 a_22300_10216 a_22212_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D37 a_3364_4822 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X739 a_33963_12403 a_33487_11828 a_33711_11850 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X740 a_35708_9001 a_37500_9006 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X741 a_32457_9520 a_32040_9564 a_32833_9564 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X742 a_36064_7612 a_35916_7168 a_35896_7612 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X743 vssd1 a_19972_9476 a_16365_5984 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X744 a_15030_7908 a_14198_8402 a_14882_8484 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X745 a_35056_10331 a_34644_10744 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X746 a_24360_9152 a_19524_11448 vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X747 a_16625_8312 a_16271_5557 vccd1 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X748 vccd1 a_21292_11351 a_21204_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X749 vssd1 a_6496_3988 a_1908_4118 vssd1 nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X750 a_3772_4032 a_3464_4076 vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X751 vccd1 a_10092_11351 a_10004_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X752 a_4069_4772 a_3949_4728 vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X753 vccd1 a_21180_4416 a_28932_4472 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X754 a_37912_12288 COMP_OUT vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X755 a_14460_11784 a_14372_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X756 vssd1 a_17696_3608 SDAC[3] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X757 a_35916_10304 a_35608_10348 vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X758 a_27748_7864 a_28428_7944 vccd1 vccd1 pfet_06v0 ad=0.2354p pd=1.95u as=0.1391p ps=1.055u w=0.535u l=0.5u
X759 vccd1 a_12244_5176 a_13216_3608 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X760 a_16814_6894 a_16694_6296 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
D38 vssd1 a_1908_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X761 a_9717_4416 a_15254_7908 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X762 a_11312_5627 a_10900_6040 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X763 a_14876_9477 a_19361_6296 a_19297_6341 vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X764 vssd1 a_3564_7864 a_1772_7864 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X765 a_22512_4476 a_22364_4032 a_22344_4476 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X766 a_21180_4416 a_27776_7124 vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
D39 a_1908_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X767 a_27880_5644 a_27328_5627 a_27676_5644 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X768 a_30488_9710 a_28040_7944 a_33172_8692 vccd1 pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X769 a_32565_12256 a_28428_7944 vssd1 vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X770 a_12780_11351 a_12692_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X771 a_15324_6608 a_21392_8392 vssd1 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X772 a_19477_5556 a_19357_6088 a_18733_6021 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X773 a_24080_6428 a_23932_6695 a_23912_6428 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X774 a_35404_10348 a_35304_10304 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X775 vssd1 a_28428_3160 SDAC[6] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X776 vssd1 a_30163_4728 a_25839_7564 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X777 a_36268_12281 a_33461_9477 a_37092_9476 vssd1 nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X778 a_27336_4476 a_25124_4472 a_26396_4032 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X779 a_32340_7908 a_29604_9880 a_32136_7908 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.1722p ps=1.24u w=0.82u l=0.6u
X780 a_29692_4076 a_27552_5176 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X781 a_20868_5556 a_20420_6087 vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X782 vssd1 a_21180_4416 a_25124_4472 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X783 a_31763_6420 a_31623_6564 a_31275_6296 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.176p ps=1.68u w=0.4u l=0.6u
X784 vssd1 a_22560_4292 a_24080_6428 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X785 a_6172_10216 a_6084_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X786 vccd1 a_27900_11351 a_27812_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D40 vssd1 a_1908_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
D41 a_2916_4822 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X787 vssd1 a_37152_5194 a_36884_6340 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X788 a_29176_7909 a_26513_7471 vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X789 vssd1 a_31677_9224 a_31797_9268 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X790 vccd1 a_22560_4292 a_33132_6744 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.3432p ps=2.44u w=0.78u l=0.5u
X791 a_1772_7864 a_3564_7864 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X792 a_22296_9180 a_20084_9176 a_21356_8736 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
D42 a_1908_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X793 a_14904_7612 a_12692_7608 a_13964_7168 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X794 vssd1 a_15383_8679 a_17241_7909 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X795 vssd1 a_29545_5904 a_29440_6044 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X796 a_15265_6040 a_12220_3205 vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X797 vssd1 a_6558_7080 a_6426_7124 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X798 a_32175_6799 a_31275_6296 vssd1 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.1224p ps=1.04u w=0.36u l=0.6u
X799 a_23980_7438 a_24435_7098 vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X800 a_10807_7909 a_3364_4822 vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X801 a_28348_11351 a_28260_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X802 a_29244_9477 a_28425_9040 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X803 vccd1 a_9408_3608 SDAC[0] vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X804 vssd1 a_2356_4118 a_20084_9176 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X805 a_27748_7864 a_28040_7944 vccd1 vccd1 pfet_06v0 ad=0.1391p pd=1.055u as=0.4268p ps=2.175u w=0.535u l=0.5u
X806 DIGITAL_OUT a_1772_7864 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X807 a_24331_11044 a_23855_11620 a_24079_11044 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X808 COMP_CLK a_33916_11000 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X809 a_25629_4728 a_23652_7608 vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X810 a_7380_5556 a_2468_4822 a_3720_5600 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4248p ps=1.94u w=1.22u l=0.5u
X811 a_25749_4772 a_25629_4728 a_25005_4728 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X812 vssd1 a_31465_5512 a_32059_4772 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X813 a_36856_7612 a_34644_7608 a_35916_7168 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X814 vccd1 a_32995_11784 a_32863_11828 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X815 a_36154_11828 a_36044_12281 a_35304_10304 vccd1 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X816 a_27648_4476 a_25536_4059 a_27336_4476 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
D43 vssd1 a_2468_4822 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X817 a_3920_4476 a_3772_4032 a_3752_4476 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X818 vccd1 a_5797_6296 a_5713_6744 vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X819 vssd1 a_33487_11828 a_33963_12403 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X820 vssd1 a_13216_3608 SDAC[1] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X821 vccd1 a_7203_6296 a_4341_6296 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X822 a_19768_7584 a_20028_7080 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X823 SC a_35708_9001 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X824 vccd1 a_4573_4728 a_4693_5348 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X825 vssd1 a_31117_7864 a_31237_7908 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X826 vccd1 a_4380_9783 a_4292_9880 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X827 vccd1 a_2356_4118 a_7652_4855 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X828 vccd1 a_2140_10216 a_2052_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X829 vssd1 a_30220_3160 a_28428_3160 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X830 vssd1 a_8157_6296 a_8277_6340 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X831 a_35896_10748 a_35056_10331 a_35608_10348 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X832 a_33912_5231 a_33511_5187 a_32855_4996 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X833 a_17850_6340 a_17730_6296 vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X834 a_35404_7212 a_27609_11448 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X835 a_22608_9180 a_20496_8763 a_22296_9180 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X836 vssd1 a_34980_6340 a_3364_4822 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
D44 a_1908_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X837 a_36268_12281 a_36084_6377 a_36884_9880 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X838 a_31561_4336 a_31144_4476 a_31937_4476 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X839 vccd1 a_22157_6088 a_22277_5556 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X840 vccd1 a_5272_6044 a_5689_5904 vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X841 a_19477_6132 a_19357_6088 a_18733_6021 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X842 a_26208_8763 a_25796_9176 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X843 vccd1 a_16252_11784 a_16164_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X844 vssd1 a_14280_9152 a_7484_5512 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X845 a_12892_3944 a_14567_4728 a_14503_4773 vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X846 vccd1 a_7068_9783 a_6980_9880 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X847 vssd1 a_21180_4416 a_21092_4472 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X848 vccd1 a_15568_5176 SDAC[2] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X849 vccd1 a_31100_9831 a_30996_9880 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
D45 a_1908_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X850 a_13653_10836 a_13533_10792 a_12909_10725 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X851 a_3464_8780 a_2912_8763 a_3260_8780 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X852 a_34174_9476 a_34054_9432 vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X853 vssd1 a_5689_5904 a_5584_6044 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X854 vccd1 a_3564_7864 a_1772_7864 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X855 a_27452_4796 a_27935_4728 a_27847_5176 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X856 vssd1 a_6496_3988 a_1908_4118 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X857 a_37500_9006 a_37108_12359 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X858 a_18376_9564 a_16576_9880 a_17436_9831 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X859 vccd1 a_17864_8648 a_17368_8692 vccd1 pfet_06v0 ad=0.4005p pd=2.12u as=0.3172p ps=1.74u w=1.22u l=0.5u
X860 a_23420_6744 a_23320_6574 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X861 a_3444_7212 a_2276_7608 a_3240_7212 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X862 a_17128_9880 a_16164_9559 a_16924_9880 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X863 a_27068_8736 a_26760_8780 vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X864 vccd1 a_12741_6341 a_13370_7908 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X865 vssd1 a_10281_4816 a_10176_4860 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X866 vccd1 a_35708_9001 SC vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X867 a_7295_4773 a_2916_4822 a_5020_6341 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X868 vssd1 a_10035_7080 a_9903_7124 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X869 vssd1 a_1772_7864 DIGITAL_OUT vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X870 vssd1 a_37196_11045 a_26163_11000 vssd1 nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
X871 COMP_CLK a_33916_11000 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X872 vssd1 a_2356_4118 a_2500_4472 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X873 vssd1 a_5129_9040 a_5024_9180 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
D46 a_2916_4822 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X874 vccd1 a_2916_4822 a_14295_5176 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X875 vssd1 a_21404_3160 a_21504_3608 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
D47 vssd1 a_1908_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X876 vccd1 a_8269_3160 a_8389_3780 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X877 vssd1 a_28428_3160 SDAC[6] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X878 vssd1 a_22803_9432 a_22671_9476 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X879 SDAC[1] a_13216_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X880 vccd1 a_11100_11784 a_11012_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X881 vccd1 a_17228_3197 a_17114_3608 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X882 a_16291_6040 a_6252_7864 vssd1 vssd1 nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
X883 a_14430_8484 a_13994_8484 a_14198_8402 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X884 a_8389_3204 a_8269_3160 a_7645_3160 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X885 vssd1 a_21180_4416 a_25796_9176 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X886 a_2912_8763 a_2500_9176 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X887 a_3668_8780 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
D48 vssd1 a_2356_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X888 DIGITAL_OUT a_1772_7864 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X889 a_11285_4773 a_10281_4816 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X890 vccd1 a_25548_11351 a_25460_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X891 vssd1 a_16926_3608 a_20420_6087 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X892 vssd1 a_37912_3205 a_34028_3160 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X893 vccd1 a_14348_11351 a_14260_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X894 vccd1 a_21871_6818 a_23927_5557 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X895 vssd1 a_22157_6088 a_22277_6132 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X896 vccd1 a_4760_6341 a_3228_3228 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X897 vssd1 a_27748_7864 a_17456_8648 vssd1 nfet_06v0 ad=0.2424p pd=1.635u as=0.341p ps=2.43u w=0.775u l=0.6u
X898 vccd1 a_4964_3608 a_6496_3988 vccd1 pfet_06v0 ad=0.367p pd=1.92u as=0.2952p ps=1.54u w=0.82u l=0.5u
X899 a_23089_9180 a_1908_4118 vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X900 a_26376_4476 a_25536_4059 a_26088_4076 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X901 a_28188_5600 a_27880_5644 vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X902 SDAC[8] a_33916_7864 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X903 a_18716_11784 a_18628_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X904 a_5129_4336 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X905 a_21180_11784 a_21092_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X906 a_22848_5176 a_22932_4728 a_22868_4772 vssd1 nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
X907 vccd1 a_27776_7124 a_21180_4416 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X908 a_2468_4822 a_27924_6340 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.4941p ps=2.03u w=1.22u l=0.5u
X909 a_1908_4118 a_6496_3988 vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X910 a_37152_5194 a_36972_7864 a_37172_4772 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X911 a_8968_7996 a_7168_8312 a_8028_8263 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X912 a_13944_7612 a_13104_7195 a_13656_7212 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X913 a_34174_10030 a_34054_9432 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X914 a_35220_4076 a_34144_9238 vccd1 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.22725p ps=1.91u w=0.505u l=0.5u
X915 a_7720_8312 a_6756_7991 a_7516_8312 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X916 a_13216_3608 a_12244_5176 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X917 vssd1 a_12244_5176 a_13216_3608 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X918 vccd1 a_2468_4822 a_6260_5176 vccd1 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X919 a_4488_7612 a_2688_7195 a_3548_7168 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
D49 a_3364_4822 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X920 vccd1 a_7292_11784 a_7204_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X921 a_35304_10304 a_36044_12281 vssd1 vssd1 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X922 vccd1 a_10527_7124 a_10983_7146 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X923 a_6060_11351 a_5972_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X924 a_3240_7212 a_2276_7608 a_3036_7212 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X925 vccd1 a_33916_11000 COMP_CLK vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X926 a_17332_9880 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X927 DIGITAL_OUT a_1772_7864 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X928 a_11548_11784 a_11460_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X929 a_3036_11351 a_2948_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X930 a_22713_9040 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X931 SDAC[3] a_17696_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X932 a_15321_7472 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X933 a_28040_7944 a_33766_10596 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X934 vccd1 a_9532_9783 a_9444_9880 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X935 a_18935_7908 a_16365_5984 a_18751_7908 vssd1 nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X936 a_5024_9180 a_2500_9176 a_4712_9180 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X937 vssd1 a_19913_4336 a_19808_4476 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X938 vssd1 a_30220_3160 a_28428_3160 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X939 a_23295_10052 a_22671_9476 a_23127_10052 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X940 vccd1 a_7884_8692 a_9408_3608 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X941 a_35896_7612 a_35056_7195 a_35608_7212 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X942 a_9308_11784 a_9220_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X943 a_14882_8484 a_14198_8402 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1656p ps=1.28u w=0.36u l=0.5u
X944 SDAC[6] a_28428_3160 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X945 vssd1 a_27776_7124 a_21180_4416 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X946 a_33916_7864 a_35708_7864 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X947 vccd1 a_4604_8215 a_4516_8312 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X948 a_22056_4076 a_21504_4059 a_21852_4076 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X949 vccd1 a_12552_9180 a_12969_9040 vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X950 vccd1 a_27935_4728 a_34980_6340 vccd1 pfet_06v0 ad=0.4941p pd=2.03u as=0.5368p ps=3.32u w=1.22u l=0.5u
X951 vccd1 a_14796_11351 a_14708_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X952 a_20495_6296 a_20196_8000 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2344p ps=1.56u w=0.82u l=0.6u
X953 vccd1 a_12580_3608 a_15568_5176 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X954 a_10035_7080 a_9385_7952 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X955 a_6679_5176 a_6133_3989 a_5020_6341 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X956 a_17676_5512 a_9717_4416 a_19655_4773 vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X957 a_8924_5127 a_8616_5176 vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X958 vccd1 a_22560_4292 a_31275_6296 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.26p ps=1.52u w=1u l=0.5u
X959 vssd1 a_23200_4728 a_22848_5176 vssd1 nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
D50 vssd1 a_1908_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X960 vssd1 a_24249_9880 a_35336_4816 vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X961 a_37152_5194 a_27856_11828 vccd1 vccd1 pfet_06v0 ad=0.4248p pd=1.94u as=0.4972p ps=3.14u w=1.13u l=0.5u
X962 a_4332_5600 a_4024_5644 vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X963 vssd1 a_23855_11620 a_24331_11044 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X964 a_32040_9564 a_29828_9559 a_31100_9831 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X965 vssd1 a_12969_9040 a_12864_9180 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X966 a_27236_6744 a_27116_6296 vccd1 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
D51 vssd1 a_2916_4822 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X967 vccd1 a_33916_7864 SDAC[8] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X968 SDAC[0] a_9408_3608 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
D52 CLK vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X969 vccd1 a_2140_11784 a_2052_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X970 vccd1 a_25374_11784 a_25242_11828 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X971 a_14540_8648 a_16325_7125 a_17904_8312 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.44955p ps=1.955u w=1.215u l=0.5u
X972 vccd1 a_37513_4416 a_36833_4476 vccd1 pfet_06v0 ad=0.3276p pd=1.62u as=0.2028p ps=1.3u w=0.78u l=0.5u
X973 a_23912_6428 a_23072_6744 a_23624_6744 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X974 vssd1 a_11123_4381 a_8479_5996 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X975 vssd1 a_15940_9880 a_17696_3608 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X976 vccd1 a_18836_7642 a_19076_11089 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X977 a_12860_7909 a_16325_7125 a_16625_8312 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X978 a_33616_4816 a_21180_4416 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X979 vssd1 a_34104_5118 a_33912_5231 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=0.2007p ps=1.475u w=0.36u l=0.6u
X980 vssd1 a_1772_7864 DIGITAL_OUT vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X981 a_3484_11351 a_3396_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X982 a_3772_8736 a_3464_8780 vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X983 a_31797_9268 a_31677_9224 a_31053_9157 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X984 a_11996_11784 a_11908_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X985 SDAC[1] a_13216_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X986 a_28129_4476 a_22560_4292 vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X987 vccd1 a_15881_4336 a_15776_4476 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X988 vccd1 a_2916_4822 a_19447_5176 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X989 a_7050_7124 a_6426_7124 a_6902_7700 vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X990 a_15324_6608 a_21392_8392 vssd1 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X991 vccd1 a_31148_11784 a_31060_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D53 vssd1 a_2916_4822 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X992 vccd1 a_11737_6384 a_11632_6428 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X993 a_9756_11784 a_9668_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X994 a_35916_10304 a_35608_10348 vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X995 a_31573_10836 a_31453_10792 a_30829_10725 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X996 a_17640_7564 a_15553_5512 vssd1 vssd1 nfet_06v0 ad=0.1248p pd=1u as=0.2112p ps=1.84u w=0.48u l=0.6u
X997 vssd1 a_35708_9001 SC vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X998 vccd1 a_7404_11351 a_7316_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X999 vssd1 a_15881_4336 a_15776_4476 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X1000 a_32352_9564 a_30240_9880 a_32040_9564 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X1001 a_9632_5556 a_9532_5512 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1002 a_15057_5557 a_15329_5996 vccd1 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1003 vssd1 a_36008_3205 a_31241_5512 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X1004 a_27776_7124 a_15324_6608 vccd1 vccd1 pfet_06v0 ad=0.2952p pd=1.54u as=0.3608p ps=2.52u w=0.82u l=0.5u
X1005 a_31465_5512 a_32404_7864 a_32340_7908 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1006 a_21891_6340 a_6252_7864 vssd1 vssd1 nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1007 a_12916_5176 a_12468_4817 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X1008 a_31750_7460 a_29739_6744 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4941p ps=2.03u w=1.22u l=0.5u
X1009 a_31750_7460 a_29739_6744 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2911p ps=1.53u w=0.82u l=0.6u
X1010 a_18836_7642 a_15553_5512 vssd1 vssd1 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X1011 a_3752_4476 a_2912_4059 a_3464_4076 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1012 a_22932_4728 a_31561_4336 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1013 a_8415_6040 a_2916_4822 a_3596_3228 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X1014 vccd1 a_17036_11351 a_16948_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1015 a_25125_4772 a_25005_4728 vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X1016 a_4693_5348 a_4573_4728 a_3949_4728 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1017 a_28425_9040 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X1018 a_23127_6040 a_20028_7080 vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1019 a_18354_6296 a_14533_5557 vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1020 a_2588_11784 a_2500_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1021 a_16365_5984 a_19972_9476 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2911p ps=1.53u w=0.82u l=0.6u
X1022 a_5724_10216 a_5636_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1023 a_9280_7996 a_7168_8312 a_8968_7996 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X1024 a_12556_4773 a_15329_5996 a_15265_6040 vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1025 a_8277_6340 a_8157_6296 a_7533_6296 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X1026 a_37649_7612 a_1908_4118 vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X1027 a_30792_9880 a_29828_9559 a_30588_9880 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1028 a_1908_4118 a_6496_3988 vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1029 a_28119_4728 a_29044_12359 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X1030 a_22277_5556 a_22157_6088 a_21533_6021 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1031 a_27847_5176 a_28527_4728 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1032 a_34364_5176 a_33912_5231 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.45p ps=2.02u w=0.78u l=0.5u
X1033 a_12741_6341 a_11737_6384 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1034 a_13994_8484 a_13370_7908 a_13826_8484 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1035 a_22000_9432 a_19361_6296 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.2344p ps=1.56u w=0.36u l=0.6u
X1036 a_22932_4728 a_31561_4336 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1037 vssd1 a_4964_3608 a_5524_3249 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1038 a_13216_3608 a_12244_5176 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1039 a_32052_5556 a_22848_5176 vccd1 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X1040 a_4828_9783 a_4740_9880 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1041 vccd1 a_21180_4416 a_26916_6040 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X1042 a_34888_9152 a_32565_12256 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X1043 a_28188_5600 a_27880_5644 vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X1044 a_36884_6340 a_36972_7864 a_35100_5996 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1045 a_1772_7864 a_3564_7864 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1046 a_21336_9180 a_20496_8763 a_21048_8780 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1047 a_37912_3205 a_22932_4728 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X1048 a_3596_3228 a_3364_4822 a_7799_5557 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1049 vccd1 a_7852_11351 a_7764_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1050 vssd1 a_21180_4416 a_34420_4472 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1051 vccd1 a_4828_11351 a_4740_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1052 COMP_CLK a_33916_11000 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1053 vccd1 a_7884_8692 a_9408_3608 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1054 SDAC[4] a_21504_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1055 SDAC[6] a_28428_3160 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1056 a_25665_6428 a_22560_4292 vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X1057 vccd1 a_23295_10052 a_23751_10030 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1058 a_2356_4118 a_13496_6366 vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1059 a_20411_6760 a_17004_3197 vccd1 vccd1 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1060 SDAC[7] a_32236_3160 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1061 a_36833_6044 a_34832_5627 a_36609_6044 vccd1 pfet_06v0 ad=0.1826p pd=1.71u as=0.1079p ps=0.935u w=0.415u l=0.5u
X1062 a_32381_11802 a_32964_10791 vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X1063 a_37513_5984 a_36609_6044 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.3276p ps=1.62u w=0.78u l=0.5u
X1064 vccd1 a_29604_9880 a_30668_7577 vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1065 vccd1 a_1772_7864 DIGITAL_OUT vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1066 a_9280_7996 a_6756_7991 a_8968_7996 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1067 vssd1 a_2468_3254 a_26241_7564 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1068 vccd1 a_17484_11351 a_17396_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1069 vccd1 a_32909_11000 a_33029_11620 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1070 a_15324_6608 a_21392_8392 vssd1 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
D54 a_1908_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1071 vccd1 a_30499_10653 a_28540_9500 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1072 vccd1 a_21180_4416 a_34420_6040 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X1073 a_1908_4118 a_6496_3988 vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.367p ps=1.92u w=1.22u l=0.5u
X1074 vssd1 a_23295_10052 a_23771_9476 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X1075 vccd1 a_36680_3205 a_35708_7864 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1076 a_12084_8312 a_2468_4822 a_9768_6574 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4248p ps=1.94u w=1.22u l=0.5u
X1077 a_8389_3780 a_8269_3160 a_7645_3160 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1078 a_9520_6744 a_9108_6423 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X1079 vccd1 a_35708_7864 a_33916_7864 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1080 vssd1 a_22560_4292 a_30352_4476 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1081 a_10281_4816 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X1082 vccd1 a_7068_10216 a_6980_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1083 a_8269_3160 a_6133_3989 vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1084 vccd1 a_15804_11784 a_15716_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1085 a_18452_4076 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
D55 a_3364_4822 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1086 vccd1 a_11324_10216 a_11236_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1087 a_30815_6341 a_29739_6744 a_30387_6744 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X1088 a_12916_5176 a_12468_4817 vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X1089 a_13029_10282 a_12909_10725 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X1090 vssd1 a_15030_7908 a_15506_7908 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X1091 vccd1 a_16365_5984 a_16271_5557 vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X1092 vssd1 a_3228_3228 a_3140_3272 vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1093 a_17128_9880 a_16576_9880 a_16924_9880 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1094 a_8820_5176 a_7652_4855 a_8616_5176 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1095 a_22277_6132 a_22157_6088 a_21533_6021 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X1096 vssd1 a_17416_6016 a_9532_5512 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X1097 vccd1 a_2356_4118 a_3060_6040 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
D56 a_1908_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1098 a_21048_8780 a_20084_9176 a_20844_8780 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1099 vccd1 a_22560_4292 a_32507_4728 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.26p ps=1.52u w=1u l=0.5u
X1100 vssd1 a_6133_8693 a_7295_4773 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1101 SDAC[1] a_13216_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1102 vccd1 a_13216_3608 SDAC[1] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1103 vccd1 a_16108_3228 a_6252_7864 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1104 a_30933_6040 a_20609_5176 vssd1 vssd1 nfet_06v0 ad=85.2f pd=0.95u as=0.3124p ps=2.3u w=0.71u l=0.6u
X1105 a_14012_4076 a_12992_3988 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X1106 a_28428_3160 a_30220_3160 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1107 vssd1 a_3564_7864 a_1772_7864 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1108 a_27131_11044 a_26655_11620 a_26879_11044 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X1109 a_20411_6760 a_6252_7864 vccd1 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X1110 a_17820_10216 a_17732_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1111 vccd1 a_25996_10747 a_25908_10791 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1112 a_3364_4822 a_34980_6340 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2911p ps=1.53u w=0.82u l=0.6u
D57 a_1908_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1113 vccd1 a_37912_3205 a_34028_3160 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1114 vccd1 a_12332_11351 a_12244_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1115 vccd1 a_2468_3254 a_10428_5870 vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1116 vccd1 a_34441_11828 a_36884_9880 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X1117 vssd1 a_23363_11000 a_23231_11044 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X1118 a_16576_9880 a_16164_9559 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1119 a_4332_5600 a_4024_5644 vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X1120 a_19797_9477 a_18793_9520 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1121 SDAC[2] a_15568_5176 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1122 vssd1 a_1908_4118 a_8176_7996 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1123 vccd1 a_27776_7124 a_21180_4416 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1124 a_33500_9006 a_28040_7944 vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1125 a_26293_6341 a_25289_6384 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1126 a_29692_4076 a_27552_5176 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X1127 a_17864_7080 a_17456_7080 a_18244_7124 vccd1 pfet_06v0 ad=0.2464p pd=2u as=0.1456p ps=1.08u w=0.56u l=0.5u
X1128 a_1772_7864 a_3564_7864 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1129 a_27048_9180 a_26208_8763 a_26760_8780 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1130 vccd1 a_29604_9880 a_32964_10791 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1131 a_4712_9180 a_2500_9176 a_3772_8736 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X1132 a_10176_4860 a_7652_4855 a_9864_4860 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1133 vccd1 a_16569_5984 a_19300_10744 vccd1 pfet_06v0 ad=0.35315p pd=1.96u as=0.2486p ps=2.01u w=0.565u l=0.5u
X1134 vssd1 a_19797_9477 a_19972_9476 vssd1 nfet_06v0 ad=0.2911p pd=1.53u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1135 a_5024_4476 a_2912_4059 a_4712_4476 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X1136 a_21852_10216 a_21764_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1137 a_11864_5644 a_11312_5627 a_11660_5644 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1138 a_34144_8693 a_30913_5557 vccd1 vccd1 pfet_06v0 ad=0.44955p pd=1.955u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1139 vccd1 a_9532_10216 a_9444_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1140 a_20732_11784 a_20644_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1141 a_8412_10216 a_8324_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1142 vssd1 a_2356_4118 a_2500_9176 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1143 SC a_35708_9001 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1144 a_9868_6744 a_9768_6574 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X1145 a_35812_7212 a_34644_7608 a_35608_7212 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1146 vccd1 a_31955_11000 a_30879_6296 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1147 a_30499_10653 a_30829_10725 a_30949_10835 vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X1148 DIGITAL_OUT a_1772_7864 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1149 SDAC[3] a_17696_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1150 vccd1 a_17696_3608 SDAC[3] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1151 a_27552_5176 a_27452_4796 vssd1 vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1152 a_13452_7212 a_13352_7168 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X1153 vssd1 a_34028_3160 a_32236_3160 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1154 vssd1 a_18836_7642 a_19076_11089 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1155 vccd1 a_26723_10216 a_26591_10260 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1156 vccd1 a_19797_9477 a_20196_8000 vccd1 pfet_06v0 ad=0.35315p pd=1.96u as=0.2486p ps=2.01u w=0.565u l=0.5u
X1157 vssd1 a_22560_4292 a_26544_4476 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1158 a_25536_4059 a_25124_4472 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X1159 a_2468_3254 a_33094_5892 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
D58 vssd1 a_1908_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1160 vccd1 a_8076_9783 a_7988_9880 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1161 a_21504_3608 a_21404_3160 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
D59 vssd1 a_1908_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1162 a_18536_10720 a_18648_4748 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X1163 a_28425_9040 a_28008_9180 a_28801_9180 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X1164 vssd1 a_27776_7124 a_21180_4416 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1165 SDAC[8] a_33916_7864 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1166 vssd1 a_33916_11000 COMP_CLK vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1167 vssd1 a_13216_3608 SDAC[1] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1168 a_37513_5984 a_36609_6044 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.14985p ps=1.145u w=0.405u l=0.6u
X1169 vccd1 a_12780_11351 a_12692_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1170 a_11304_8780 a_10752_8763 a_11100_8780 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1171 a_25289_6384 a_22560_4292 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X1172 vssd1 a_13529_5904 a_13424_6044 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X1173 a_30028_11351 a_29940_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1174 vccd1 a_14616_9477 a_12188_7864 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1175 a_35677_5644 a_34420_6040 a_35424_5644 vccd1 pfet_06v0 ad=0.101p pd=0.905u as=0.19315p ps=1.27u w=0.505u l=0.5u
X1176 vccd1 a_27215_10260 a_27671_10282 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
D60 a_2468_3254 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1177 vccd1 a_6844_11784 a_6756_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1178 vccd1 a_13496_6366 a_2356_4118 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1179 a_5612_11351 a_5524_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1180 a_29896_4076 a_28932_4472 a_29692_4076 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1181 vccd1 a_33916_11000 COMP_CLK vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1182 a_32352_9564 a_29828_9559 a_32040_9564 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1183 a_22260_4076 a_21092_4472 a_22056_4076 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1184 a_25184_6428 a_23072_6744 a_24872_6428 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X1185 SDAC[7] a_32236_3160 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1186 a_27336_4476 a_25536_4059 a_26396_4032 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1187 vccd1 a_37500_4728 a_37396_5176 vccd1 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1188 a_21871_5250 a_6252_7864 vccd1 vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X1189 a_12068_5644 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X1190 a_26088_4076 a_25124_4472 a_25884_4076 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1191 vccd1 a_4229_3160 a_4145_3608 vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1192 a_8086_7700 a_7254_7124 a_7918_7700 vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1193 a_24540_9783 a_24452_9880 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1194 a_18760_8692 a_18828_9199 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1195 a_1908_4118 a_6496_3988 vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1196 a_12600_7909 a_12860_7909 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X1197 a_6902_7700 a_6426_7124 vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1198 a_11632_6428 a_9108_6423 a_11320_6428 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1199 a_15244_11351 a_15156_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1200 vccd1 a_28348_11351 a_28260_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1201 vccd1 a_23196_10216 a_23108_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1202 vssd1 a_6496_3988 a_1908_4118 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1203 a_37172_4772 a_27856_11828 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1204 vccd1 a_9980_10216 a_9892_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1205 a_34144_8693 a_31465_5512 a_34144_9238 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1206 vssd1 a_16364_6296 a_14567_4728 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1207 vssd1 a_4905_7472 a_4800_7612 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X1208 a_13656_7212 a_12692_7608 a_13452_7212 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1209 a_8860_10216 a_8772_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1210 a_29545_5904 a_22560_4292 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
D61 a_1908_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1211 a_7516_8312 a_7416_8142 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1212 a_36064_10748 a_35916_10304 a_35896_10748 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1213 a_3668_4076 a_2500_4472 a_3464_4076 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1214 a_7740_11784 a_7652_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1215 a_37500_9006 a_37108_12359 vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X1216 vssd1 a_33461_9477 a_37780_9568 vssd1 nfet_06v0 ad=0.2344p pd=1.56u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1217 vccd1 a_33724_9432 a_30471_6296 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1218 vccd1 a_2356_4118 a_10340_9176 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X1219 a_28055_4773 a_27935_4728 vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1220 a_7526_7700 a_7050_7124 a_7254_7124 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X1221 vssd1 a_6133_8693 a_6140_4728 vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1222 vssd1 a_32909_11000 a_33029_11044 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1223 vssd1 a_17696_3608 SDAC[3] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1224 vssd1 a_35708_9001 SC vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1225 a_10787_8312 a_3364_4822 a_10599_8312 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1226 vccd1 a_13216_3608 SDAC[1] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1227 a_36680_3205 a_30981_5996 vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X1228 a_16364_6296 a_16694_6296 a_16814_6894 vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1229 a_19768_7584 a_20028_7080 vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X1230 a_36856_7612 a_35056_7195 a_35916_7168 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1231 a_27116_6296 a_26804_7953 vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X1232 a_30476_11351 a_30388_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1233 a_35608_7212 a_34644_7608 a_35404_7212 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1234 vccd1 a_36008_3205 a_31241_5512 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1235 vssd1 a_28428_3160 SDAC[6] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1236 vccd1 a_33766_10596 a_28040_7944 vccd1 pfet_06v0 ad=0.4941p pd=2.03u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1237 a_21180_4416 a_27776_7124 vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1238 vccd1 a_20096_10688 a_18940_7080 vccd1 pfet_06v0 ad=0.35315p pd=1.96u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1239 vccd1 a_34980_6340 a_3364_4822 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1240 vssd1 a_13533_10792 a_13653_10836 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1241 vccd1 a_18793_9520 a_18688_9564 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
D62 vssd1 a_2468_3254 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1242 a_1692_10216 a_1604_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1243 a_17372_11784 a_17284_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1244 vssd1 a_21504_3608 SDAC[4] vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1245 a_33407_5231 a_32507_4728 vssd1 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.1224p ps=1.04u w=0.36u l=0.6u
X1246 a_7799_5557 a_8479_5996 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1247 vccd1 a_29804_10216 a_29716_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1248 vccd1 a_22524_11784 a_22436_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1249 a_35230_10052 a_35090_9432 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1656p ps=1.28u w=0.36u l=0.5u
X1250 a_35668_4476 a_34832_4059 a_35424_4076 vssd1 nfet_06v0 ad=62.1f pd=0.705u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1251 a_9653_4472 a_2468_3254 vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1252 a_17696_3608 a_15940_9880 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1253 a_14911_4773 a_2916_4822 a_12892_3944 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X1254 a_34069_6040 a_28040_7944 vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1255 a_12077_4520 a_11285_4773 vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1256 a_30949_10282 a_30829_10725 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X1257 vssd1 a_32236_3160 SDAC[7] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1258 a_26556_8780 a_26456_8736 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X1259 a_23304_4476 a_21504_4059 a_22364_4032 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1260 a_12580_3608 a_12132_3249 vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
D63 a_2356_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1261 a_15692_11351 a_15604_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1262 a_27653_10052 a_27533_9432 a_26909_9432 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1263 a_36833_6044 a_34420_6040 a_36609_6044 vssd1 nfet_06v0 ad=0.2898p pd=2.33u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1264 a_30723_9085 a_31053_9157 a_31173_8714 vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1265 a_24872_6428 a_23072_6744 a_23932_6695 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1266 vccd1 a_1692_7080 a_1604_7124 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1267 vssd1 a_21392_8392 a_15324_6608 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X1268 a_18248_4076 a_17696_4059 a_18044_4076 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1269 vssd1 a_8479_5996 a_8415_6040 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1270 vssd1 a_28040_7944 a_29075_6875 vssd1 nfet_06v0 ad=0.2288p pd=1.58u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1271 a_33487_11828 a_32863_11828 a_33319_11828 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1272 a_6496_3988 a_4964_3608 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1273 a_3260_4076 a_3160_4032 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X1274 a_26768_5176 a_19052_8648 a_26564_5176 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1275 vccd1 a_25374_11784 a_37108_12359 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
D64 a_2356_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1276 vssd1 a_26655_11620 a_27131_11044 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X1277 a_32855_4996 a_33511_5187 a_33407_5231 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.1313p ps=1.025u w=0.505u l=0.5u
X1278 a_3932_9783 a_3844_9880 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1279 a_24540_10216 a_24452_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1280 vssd1 a_22560_4292 a_31763_6420 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=0.134p ps=1.1u w=0.36u l=0.6u
X1281 a_2356_4118 a_13496_6366 vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1282 vssd1 a_25629_4728 a_25749_4772 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1283 a_30996_9880 a_29828_9559 a_30792_9880 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1284 a_23420_11784 a_23332_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1285 vssd1 a_25866_11828 a_26342_12404 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1286 a_21504_3608 a_21404_3160 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1287 a_15776_4476 a_13252_4472 a_15464_4476 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1288 a_2912_4059 a_2500_4472 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X1289 a_19089_6744 a_16365_5984 a_14876_9477 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1290 vccd1 a_21404_3160 a_21504_3608 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1291 a_32872_6686 a_32384_6384 a_33132_6744 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1292 a_8269_3160 a_6133_3989 vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1293 a_12172_5600 a_11864_5644 vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X1294 a_30778_7124 a_30668_7577 vccd1 vccd1 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1295 SC a_35708_9001 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1296 SDAC[1] a_13216_3608 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1297 vssd1 a_13216_3608 SDAC[1] vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1298 a_18388_4728 a_17640_7564 a_19028_5308 vccd1 pfet_06v0 ad=0.2464p pd=2u as=0.1736p ps=1.18u w=0.56u l=0.5u
X1299 vccd1 CLK a_21392_8392 vccd1 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X1300 a_7799_5557 a_5797_6296 a_3596_3228 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1301 vssd1 a_36268_12281 a_35304_10304 vssd1 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X1302 a_30352_4476 a_30204_4032 a_30184_4476 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1303 vccd1 a_22972_11784 a_22884_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1304 vccd1 a_14524_4032 a_14420_4076 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1305 a_1692_5079 a_1604_5176 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D65 vssd1 a_2468_3254 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1306 a_21740_11351 a_21652_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1307 a_13352_7168 a_17456_7080 a_17368_7124 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1308 a_10540_11351 a_10452_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1309 a_31117_4728 a_23599_5996 vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1310 vssd1 a_22560_4292 a_36064_10748 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1311 a_11123_4381 a_11453_4453 a_11573_4010 vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1312 vssd1 a_19052_8648 a_26513_7471 vssd1 nfet_06v0 ad=0.1209p pd=0.985u as=0.1209p ps=0.985u w=0.465u l=0.6u
X1313 a_15506_7908 a_15030_7908 a_15254_7908 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X1314 a_8300_11351 a_8212_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1315 vccd1 a_15324_6608 a_13496_6366 vccd1 pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X1316 a_33724_9432 a_34054_9432 a_34174_10030 vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1317 vssd1 a_15940_9880 a_17696_3608 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1318 a_33912_5231 a_33616_4816 a_32855_4996 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.25375p ps=1.51u w=0.505u l=0.5u
X1319 a_13572_5176 a_12916_5176 vccd1 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X1320 a_3596_3228 a_5797_6296 a_8007_6040 vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1321 vssd1 a_1908_4118 a_21504_9180 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1322 a_32236_3160 a_34028_3160 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1323 a_12077_4520 a_11285_4773 vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1324 a_17456_7080 a_17456_8648 vccd1 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X1325 vssd1 a_18354_6296 a_18474_6340 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1326 vccd1 a_26356_10260 a_34980_3249 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1327 a_13846_7908 a_13370_7908 vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1328 a_30588_9880 a_30488_9710 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1329 vccd1 a_33616_4816 a_33511_5187 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X1330 a_36084_6377 a_32381_11802 vssd1 vssd1 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X1331 a_31465_5512 a_28040_7944 vccd1 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X1332 vccd1 a_19164_11784 a_19076_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1333 a_29132_11351 a_29044_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1334 a_17904_8312 a_11285_4773 vccd1 vccd1 pfet_06v0 ad=0.44955p pd=1.955u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1335 vccd1 a_12244_5176 a_13216_3608 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1336 vssd1 a_30879_6296 a_30815_6341 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1337 a_7156_6040 a_5713_6744 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1338 a_19089_6744 a_19361_6296 vccd1 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1339 a_23444_7608 a_23756_7080 a_23652_7608 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1340 a_25698_11828 a_25242_11828 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1341 a_30499_10653 a_30829_10725 a_30949_10282 vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1342 vccd1 a_37500_9006 a_35708_9001 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
D66 a_2468_4822 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1343 vssd1 a_13496_6366 a_2356_4118 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1344 a_15216_7612 a_12692_7608 a_14904_7612 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1345 vccd1 a_6060_11351 a_5972_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1346 a_8176_7996 a_8028_8263 a_8008_7996 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1347 vssd1 a_1772_7864 DIGITAL_OUT vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1348 vccd1 a_3036_11351 a_2948_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1349 SDAC[3] a_17696_3608 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1350 a_21871_6818 a_6252_7864 vccd1 vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X1351 a_35737_4428 a_35424_4076 vccd1 vccd1 pfet_06v0 ad=0.1521p pd=1.105u as=0.3975p ps=2.185u w=0.585u l=0.5u
X1352 vssd1 a_29512_4773 a_22803_9432 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X1353 vssd1 a_21504_3608 SDAC[4] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1354 a_9768_6574 a_2468_4822 a_11860_7908 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1355 a_29772_4773 a_24809_11448 a_32977_3989 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
D67 a_2356_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1356 a_9864_4860 a_7652_4855 a_8924_5127 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X1357 a_21180_4416 a_27776_7124 vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
D68 vssd1 a_1908_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1358 a_24135_6040 a_20868_5556 vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1359 vccd1 a_10428_5870 a_7416_8142 vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X1360 vssd1 a_35708_7864 a_33916_7864 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1361 vccd1 a_6440_9152 a_3564_7864 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1362 a_7720_8312 a_7168_8312 a_7516_8312 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1363 vssd1 a_37513_5984 a_37465_6040 vssd1 nfet_06v0 ad=0.14985p pd=1.145u as=48.6f ps=0.645u w=0.405u l=0.6u
X1364 a_29356_10216 a_29268_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1365 a_2588_9783 a_2500_9880 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1366 a_33768_7608 a_33096_7124 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X1367 a_33768_7124 a_33096_7124 vccd1 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4005p ps=2.12u w=1.22u l=0.5u
X1368 a_3444_7212 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X1369 a_6148_7908 a_4257_6744 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1370 a_20063_4773 a_2916_4822 a_17676_5512 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X1371 vccd1 a_3619_4728 a_3160_4032 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1372 a_4380_10216 a_4292_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1373 a_26241_7564 a_26513_7471 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.2288p ps=1.58u w=0.36u l=0.6u
X1374 a_27776_7124 a_15324_6608 vccd1 vccd1 pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X1375 vssd1 a_21392_8392 a_15324_6608 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X1376 a_31144_4476 a_28932_4472 a_30204_4032 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X1377 vccd1 a_14012_11784 a_13924_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D69 vssd1 a_2356_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1378 vccd1 a_32404_7864 a_33500_9006 vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1379 a_36008_3205 a_35428_3608 vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X1380 a_23052_7564 a_3364_4822 a_25159_7125 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1381 a_5797_6296 a_8310_7146 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X1382 vssd1 a_26723_10216 a_26591_10260 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X1383 vccd1 a_17640_7564 a_21871_5250 vccd1 pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
X1384 a_7884_8692 a_7428_9176 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2344p ps=1.56u w=0.82u l=0.6u
X1385 a_29580_11351 a_29492_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1386 a_18380_11351 a_18292_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1387 a_1692_8648 a_1604_8692 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1388 a_30387_6744 a_30471_6296 a_30407_6341 vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1389 vccd1 a_15940_9880 a_17696_3608 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1390 a_29344_4059 a_28932_4472 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
D70 a_2468_4822 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1391 a_14112_7612 a_13964_7168 a_13944_7612 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1392 a_18648_4748 a_18940_7080 a_20832_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X1393 vssd1 a_25374_11784 a_37108_12359 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1394 vssd1 a_31453_10792 a_31573_10836 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1395 vccd1 a_3484_11351 a_3396_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1396 a_17436_9831 a_17128_9880 vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X1397 vccd1 a_2356_4118 a_13252_4472 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
D71 a_16108_3228 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1398 vccd1 a_29804_11784 a_29716_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1399 a_27533_9432 a_26293_6341 vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1400 SDAC[1] a_13216_3608 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1401 a_20028_7080 a_19052_8648 vssd1 vssd1 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X1402 vccd1 a_32380_5870 a_31509_7864 vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X1403 a_7924_8312 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X1404 vccd1 a_5689_5904 a_5584_6044 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X1405 a_21203_7517 a_21533_7589 a_21653_7146 vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1406 a_28119_4728 a_29044_12359 vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X1407 a_34678_9698 a_35090_9432 a_35230_10052 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1408 a_7918_7700 a_7254_7124 vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1409 vccd1 a_22803_9432 a_22671_9476 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1410 a_18768_5308 a_18648_4748 vccd1 vccd1 pfet_06v0 ad=0.224p pd=1.36u as=0.389p ps=2.02u w=0.56u l=0.5u
X1411 a_4828_11784 a_4740_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1412 a_31677_9224 a_22932_4728 vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
D72 vssd1 a_2468_4822 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1413 a_1772_7864 a_3564_7864 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1414 vccd1 a_24675_4728 a_23320_6574 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1415 vccd1 a_13496_6366 a_2356_4118 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1416 vssd1 a_25996_10747 a_25908_10791 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1417 vccd1 CLK a_21392_8392 vccd1 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X1418 a_31456_4476 a_29344_4059 a_31144_4476 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
D73 a_1908_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1419 a_10599_8312 a_11279_7864 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1420 a_19913_4336 a_19496_4476 a_20289_4476 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X1421 a_18244_8692 a_16365_5984 vccd1 vccd1 pfet_06v0 ad=0.1456p pd=1.08u as=0.4005p ps=2.12u w=0.56u l=0.5u
X1422 a_19656_7909 a_19916_7909 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X1423 vssd1 a_2356_4118 a_16164_9559 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1424 a_9761_7996 a_1908_4118 vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
D74 a_2916_4822 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1425 a_16512_9120 a_16325_7125 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.2344p ps=1.56u w=0.36u l=0.6u
X1426 vssd1 a_17228_3197 a_16926_3608 vssd1 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X1427 a_14012_4076 a_12992_3988 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1428 a_27935_4728 a_30668_7577 vssd1 vssd1 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X1429 vccd1 a_5129_9040 a_5024_9180 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X1430 a_17576_9176 a_17456_8648 vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1431 a_5281_7612 a_1908_4118 vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X1432 vccd1 a_14460_11784 a_14372_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1433 vccd1 a_15553_5512 a_17640_7564 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1434 a_36044_12281 a_32481_11846 vssd1 vssd1 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X1435 vccd1 a_6133_8693 a_7428_9176 vccd1 pfet_06v0 ad=0.35315p pd=1.96u as=0.2486p ps=2.01u w=0.565u l=0.5u
X1436 a_26760_8780 a_25796_9176 a_26556_8780 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1437 vccd1 a_27336_4476 a_27753_4336 vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X1438 vssd1 a_35737_4428 a_35668_4476 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=62.1f ps=0.705u w=0.36u l=0.6u
X1439 vccd1 a_2356_4118 a_10900_6040 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X1440 a_15324_6608 a_21392_8392 vssd1 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X1441 a_32236_3160 a_34028_3160 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1442 vssd1 a_26163_11000 a_26031_11044 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X1443 vccd1 a_11285_4773 a_11796_4817 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1444 a_27676_5644 a_27236_6340 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X1445 a_15673_6040 a_15553_5512 a_12556_4773 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X1446 a_5129_9040 a_4712_9180 a_5505_9180 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X1447 vssd1 a_33916_7864 SDAC[8] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1448 a_17228_3197 a_20495_6296 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1449 a_31080_9564 a_30240_9880 a_30792_9880 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1450 vccd1 a_27068_8736 a_26964_8780 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1451 vssd1 a_1908_4118 a_36064_7612 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1452 vccd1 a_35708_7864 a_33916_7864 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1453 vccd1 a_18376_9564 a_18793_9520 vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X1454 vccd1 a_25866_11828 a_26302_11828 vccd1 pfet_06v0 ad=0.1656p pd=1.28u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1455 a_32136_7908 a_28040_7944 vssd1 vssd1 nfet_06v0 ad=0.1722p pd=1.24u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1456 a_31248_9564 a_31100_9831 a_31080_9564 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1457 vccd1 a_28757_3989 a_29044_12359 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1458 a_3619_4728 a_3949_4728 a_4069_4772 vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X1459 a_7156_6040 a_7484_5512 a_3720_5600 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1460 vccd1 a_22748_10216 a_22660_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1461 a_33094_5892 a_31465_5512 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2911p ps=1.53u w=0.82u l=0.6u
X1462 a_35100_5996 a_36972_7864 a_37092_6744 vccd1 pfet_06v0 ad=0.4248p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1463 a_6133_3989 a_5129_4336 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1464 a_30549_5557 a_29545_5904 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1465 a_10428_10216 a_10340_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1466 a_25374_11784 a_37513_5984 vccd1 vccd1 pfet_06v0 ad=0.6561p pd=3.51u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1467 SDAC[8] a_33916_7864 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1468 a_23127_10052 a_22671_9476 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1469 a_34832_4059 a_34420_4472 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1470 a_36884_8312 a_28169_10260 a_26163_11000 vccd1 pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1471 a_10528_6428 a_10380_6695 a_10360_6428 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1472 a_31173_8714 a_31053_9157 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X1473 a_14524_4032 a_14216_4076 vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X1474 a_16576_9880 a_16164_9559 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X1475 SDAC[4] a_21504_3608 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1476 vssd1 a_21504_3608 SDAC[4] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1477 vccd1 a_37912_12288 a_16108_3228 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1478 a_10380_6695 a_10072_6744 vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
D75 vssd1 a_2356_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1479 a_33943_11850 a_33487_11828 a_33711_11850 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X1480 vssd1 a_37500_9006 a_35708_9001 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1481 vccd1 a_16512_9120 a_15553_5512 vccd1 pfet_06v0 ad=0.35315p pd=1.96u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1482 a_21392_8392 CLK vccd1 vccd1 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X1483 a_23363_11000 a_37513_4416 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1484 vssd1 a_32236_3160 SDAC[7] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1485 vccd1 a_6252_7864 a_20609_5176 vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1486 vssd1 a_19768_7584 a_18236_7864 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X1487 a_13452_7212 a_13352_7168 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1488 a_6133_3989 a_5129_4336 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1489 a_6148_7908 a_2468_3254 a_2936_7168 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1490 vccd1 a_20495_6296 a_20922_3608 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4087p ps=1.89u w=1.22u l=0.5u
X1491 a_30549_5557 a_29545_5904 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1492 vccd1 a_35737_5996 a_35677_5644 vccd1 pfet_06v0 ad=0.3975p pd=2.185u as=0.101p ps=0.905u w=0.505u l=0.5u
X1493 vccd1 a_37152_5194 a_35100_5996 vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X1494 vssd1 a_2356_4118 a_10340_9176 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1495 a_15483_8723 a_15383_8679 vccd1 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.4334p ps=2.85u w=0.985u l=0.5u
X1496 a_9633_4006 a_9717_4416 a_9653_4472 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1497 vssd1 a_21392_8392 a_15324_6608 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X1498 vssd1 a_14975_4728 a_14911_4773 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1499 vccd1 a_27776_7124 a_21180_4416 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1500 a_26754_11828 a_26070_11828 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1656p ps=1.28u w=0.36u l=0.5u
X1501 vccd1 a_24809_11448 a_34292_8648 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1502 a_10657_4860 a_1908_4118 vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X1503 a_16325_7125 a_15321_7472 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1504 a_23707_11044 a_23231_11044 vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1505 a_37435_3204 a_28119_4728 a_32380_5870 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1506 a_16924_11784 a_16836_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1507 SDAC[3] a_17696_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1508 a_24675_4728 a_25005_4728 a_25125_4772 vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X1509 vccd1 a_9084_9783 a_8996_9880 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1510 vccd1 a_3772_8736 a_3668_8780 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1511 vccd1 a_23304_4476 a_23721_4336 vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X1512 a_14524_4032 a_14216_4076 vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X1513 a_35737_5996 a_35424_5644 vccd1 vccd1 pfet_06v0 ad=0.1521p pd=1.105u as=0.3975p ps=2.185u w=0.585u l=0.5u
X1514 vssd1 a_37196_11045 a_37108_11089 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1515 a_30184_4476 a_29344_4059 a_29896_4076 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1516 vccd1 a_23200_4728 a_22660_5176 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X1517 a_23147_9476 a_22671_9476 vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1518 a_6372_8312 a_6252_7864 a_2936_7168 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4248p ps=1.94u w=1.22u l=0.5u
X1519 vccd1 a_17456_8648 a_18828_9199 vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1520 vssd1 a_34678_9698 a_34818_9476 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1521 a_23624_6744 a_23072_6744 a_23420_6744 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1522 a_26723_10216 a_37273_7472 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1523 a_11573_4010 a_11453_4453 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X1524 a_10876_10216 a_10788_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1525 vssd1 a_16108_3228 a_18388_4728 vssd1 nfet_06v0 ad=0.104p pd=0.92u as=0.14p ps=1.1u w=0.4u l=0.6u
X1526 vccd1 a_31677_9224 a_31797_8692 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1527 SDAC[1] a_13216_3608 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1528 a_24249_9880 a_23519_9476 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X1529 a_3820_5644 a_3720_5600 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X1530 vccd1 a_12220_3205 a_12132_3249 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1531 COMP_CLK a_33916_11000 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1532 a_21504_9180 a_21356_8736 a_21336_9180 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1533 a_18474_6340 a_18354_6296 a_17730_6296 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X1534 vssd1 a_2468_3254 a_11003_9476 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1535 vccd1 a_23721_4336 a_23616_4476 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X1536 a_36609_6044 a_34832_5627 a_35737_5996 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1989p ps=1.465u w=0.36u l=0.6u
X1537 a_3364_4822 a_34980_6340 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.4941p ps=2.03u w=1.22u l=0.5u
X1538 vccd1 a_33916_7864 SDAC[8] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1539 a_13029_10835 a_12909_10725 vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X1540 a_32833_9564 a_22560_4292 vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X1541 a_27047_10260 a_26591_10260 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1542 a_6440_9152 a_5909_7125 vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X1543 SDAC[4] a_21504_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1544 vccd1 a_17640_7564 a_21871_6818 vccd1 pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
X1545 vssd1 a_23721_4336 a_23616_4476 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X1546 vccd1 a_19913_4336 a_19808_4476 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X1547 a_35424_4076 a_34420_4472 a_35220_4076 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1548 vssd1 a_36680_3205 a_35708_7864 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X1549 vccd1 a_10380_6695 a_10276_6744 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1550 vccd1 a_12077_4520 a_12197_3988 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1551 SDAC[7] a_32236_3160 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1552 a_25367_7608 a_3364_4822 vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1553 a_9520_6744 a_9108_6423 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1554 a_14295_5176 a_14567_4728 a_12892_3944 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1555 a_20615_6340 a_20495_6296 a_20431_6340 vssd1 nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1556 a_28348_11784 a_28260_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1557 vccd1 a_2588_10216 a_2500_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1558 a_15324_6608 a_21392_8392 vssd1 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X1559 a_2688_7195 a_2276_7608 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
D76 vssd1 a_2468_4822 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1560 a_1908_4118 a_6496_3988 vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1561 a_29075_6875 a_26456_8736 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1562 a_23828_6744 a_22560_4292 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X1563 vssd1 a_4964_3608 a_6496_3988 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1564 a_26088_4076 a_25536_4059 a_25884_4076 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1565 vccd1 a_33487_11828 a_33943_11850 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1566 a_22157_7656 a_20495_6296 vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1567 a_16924_9880 a_16824_9710 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X1568 a_37465_6040 a_22560_4292 a_36833_6044 vssd1 nfet_06v0 ad=48.6f pd=0.645u as=0.3123p ps=2.38u w=0.405u l=0.6u
X1569 vssd1 a_6133_8693 a_7428_9176 vssd1 nfet_06v0 ad=0.2344p pd=1.56u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1570 a_32507_4728 a_32855_4996 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X1571 vssd1 a_13496_6366 a_2356_4118 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1572 SDAC[3] a_17696_3608 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1573 a_24976_3608 a_24876_3160 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1574 a_30163_4728 a_30493_4728 a_30613_4772 vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X1575 a_21048_8780 a_20496_8763 a_20844_8780 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1576 a_23927_5557 a_17640_7564 a_24115_5557 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1577 a_32384_6384 a_21180_4416 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X1578 a_1692_11351 a_1604_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1579 a_21504_3608 a_21404_3160 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1580 vssd1 a_5972_3608 a_25312_5556 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1581 a_29244_9477 a_28425_9040 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1582 a_18536_10720 a_18648_4748 vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X1583 vccd1 a_33500_9006 a_30488_9710 vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X1584 a_30913_5557 a_30981_5996 a_30933_6040 vssd1 nfet_06v0 ad=0.21175p pd=1.41u as=85.2f ps=0.95u w=0.71u l=0.6u
X1585 a_3260_4076 a_3160_4032 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1586 a_37904_7864 a_26723_10216 vccd1 vccd1 pfet_06v0 ad=0.2486p pd=2.01u as=0.35315p ps=1.96u w=0.565u l=0.5u
X1587 vccd1 a_18716_11784 a_18628_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1588 vccd1 a_28460_10216 a_28372_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1589 a_10428_5870 a_10871_7864 vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1590 vccd1 a_13216_3608 SDAC[1] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1591 vccd1 a_21180_11784 a_21092_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1592 vccd1 a_2468_3254 a_13900_4728 vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1593 vccd1 a_37273_10608 a_37168_10748 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X1594 a_1692_9783 a_1604_9880 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1595 a_28320_9180 a_25796_9176 a_28008_9180 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1596 vccd1 a_30028_11351 a_29940_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1597 a_27856_11828 a_27126_11850 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X1598 vccd1 a_5612_11351 a_5524_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1599 a_22289_4772 a_19052_8648 a_22085_4772 vssd1 nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1600 vccd1 a_18388_4728 a_15329_5996 vccd1 pfet_06v0 ad=0.389p pd=2.02u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1601 a_26513_7471 a_17228_3197 vssd1 vssd1 nfet_06v0 ad=0.1209p pd=0.985u as=0.2046p ps=1.81u w=0.465u l=0.6u
X1602 a_33461_9477 a_32457_9520 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1603 a_17696_3608 a_15940_9880 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1604 a_13533_10792 a_10787_8312 vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1605 vccd1 a_36856_7612 a_37273_7472 vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X1606 vssd1 a_12077_4520 a_12197_4564 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1607 a_21653_7146 a_21533_7589 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X1608 vssd1 a_16512_9120 a_15553_5512 vssd1 nfet_06v0 ad=0.2344p pd=1.56u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1609 a_19361_6296 a_19913_4336 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1610 a_20629_4772 a_19524_11448 vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1611 a_28908_10216 a_28820_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1612 vccd1 a_11548_11784 a_11460_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1613 vssd1 a_12741_6341 a_13370_7908 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X1614 vccd1 a_15244_11351 a_15156_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1615 vssd1 a_21392_8392 a_15324_6608 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X1616 a_14280_9152 a_14540_8648 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X1617 a_3932_10216 a_3844_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1618 a_27880_5644 a_26916_6040 a_27676_5644 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1619 a_12741_6341 a_11737_6384 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1620 a_19612_11784 a_19524_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1621 vccd1 a_9308_11784 a_9220_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1622 a_27215_10260 a_26591_10260 a_27047_10260 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1623 a_30252_11784 a_30164_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1624 vssd1 a_33724_9432 a_30471_6296 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1625 a_26292_4076 a_22560_4292 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X1626 vccd1 a_28188_5600 a_28084_5644 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1627 a_11320_6428 a_9108_6423 a_10380_6695 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
D77 vssd1 a_2356_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1628 a_5020_6341 a_3364_4822 a_6679_5176 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
D78 vssd1 a_2468_3254 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1629 a_23652_7124 a_23107_5557 vccd1 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X1630 a_23652_7608 a_23107_5557 a_23444_7608 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1631 a_22157_7656 a_20495_6296 vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1632 vccd1 a_17696_3608 SDAC[3] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1633 vssd1 a_24876_3160 a_24976_3608 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1634 a_17932_11351 a_17844_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1635 vccd1 a_27776_7124 a_21180_4416 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1636 vccd1 a_37904_7864 a_28428_7944 vccd1 pfet_06v0 ad=0.35315p pd=1.96u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1637 a_16689_6040 a_16569_5984 a_16485_6040 vssd1 nfet_06v0 ad=0.1517p pd=1.19u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1638 a_24311_11598 a_23855_11620 a_24079_11044 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X1639 vccd1 a_30476_11351 a_30388_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1640 SDAC[4] a_21504_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1641 a_22560_4292 a_25312_5556 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1642 a_11860_7908 a_9633_4006 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1643 a_32381_11802 a_32964_10791 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X1644 a_4573_4728 a_4965_4728 vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1645 a_31226_7124 a_28040_7944 a_27935_4728 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3477p ps=1.79u w=1.22u l=0.5u
X1646 a_32565_12256 a_28428_7944 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1647 a_8188_11784 a_8100_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1648 vccd1 a_27533_9432 a_27653_10052 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1649 a_12444_11784 a_12356_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1650 a_29604_9880 a_29156_9521 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X1651 a_36833_4476 a_22560_4292 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X1652 vccd1 a_21504_3608 SDAC[4] vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1653 a_5689_5904 a_5272_6044 a_6065_6044 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X1654 vssd1 a_37273_10608 a_37168_10748 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X1655 a_32995_11784 a_37273_10608 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1656 a_32059_4772 a_30471_6296 a_27564_6296 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1657 a_12600_7909 a_12860_7909 vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X1658 a_17696_3608 a_15940_9880 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1659 a_15057_5557 a_15737_5996 a_12556_4773 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
D79 vssd1 a_1908_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1660 vccd1 a_32565_12256 a_32481_11846 vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1661 a_15324_6608 a_21392_8392 vssd1 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.2134p ps=1.85u w=0.485u l=0.6u
X1662 SDAC[7] a_32236_3160 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
D80 a_2468_4822 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1663 a_15881_4336 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X1664 a_32932_7908 a_29604_9880 a_32748_7908 vssd1 nfet_06v0 ad=0.1148p pd=1.1u as=0.1312p ps=1.14u w=0.82u l=0.6u
X1665 a_5612_9783 a_5524_9880 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1666 a_20922_3608 a_19052_8648 a_20028_7080 vccd1 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
D81 a_2468_3254 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1667 vccd1 a_11996_11784 a_11908_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1668 vccd1 a_15324_6608 a_13496_6366 vccd1 pfet_06v0 ad=0.3608p pd=2.52u as=0.2952p ps=1.54u w=0.82u l=0.5u
X1669 vccd1 a_15692_11351 a_15604_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1670 a_31955_11000 a_32285_11000 a_32405_11598 vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1671 a_19447_5176 a_9717_4416 a_17676_5512 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1672 a_11632_6428 a_9520_6744 a_11320_6428 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X1673 vccd1 a_9756_11784 a_9668_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1674 a_1908_4118 a_6496_3988 vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1675 vssd1 a_27776_7124 a_21180_4416 vssd1 nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1676 vssd1 a_1908_4118 a_3920_9180 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1677 a_23535_6040 a_20411_6760 a_23107_5557 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X1678 a_26513_7471 a_17640_7564 a_26768_5176 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1679 a_4024_5644 a_3060_6040 a_3820_5644 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1680 vccd1 a_5276_10216 a_5188_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1681 vssd1 a_15737_5996 a_15673_6040 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1682 vssd1 a_21180_4416 a_28932_4472 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1683 a_32909_11000 a_24607_5996 vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1684 a_20832_10260 a_16365_5984 vccd1 vccd1 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1685 a_30949_10835 a_30829_10725 vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X1686 a_16833_7909 a_11279_7864 vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1687 vccd1 a_14280_9152 a_7484_5512 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1688 a_15697_7612 a_1908_4118 vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X1689 a_19052_8648 a_19300_10744 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.35315p ps=1.96u w=1.22u l=0.5u
X1690 a_3036_11784 a_2948_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1691 vssd1 a_27533_9432 a_27653_9476 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1692 a_22260_4076 a_22560_4292 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X1693 vssd1 a_7050_7124 a_7526_7700 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
D82 a_2356_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1694 a_21504_3608 a_21404_3160 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1695 vssd1 a_25312_5556 a_22560_4292 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1696 a_15324_6608 a_21392_8392 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1697 vccd1 a_13216_3608 SDAC[1] vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1698 a_3464_8780 a_2500_9176 a_3260_8780 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1699 a_4380_11351 a_4292_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1700 a_21392_8392 CLK vccd1 vccd1 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X1701 vccd1 a_2588_11784 a_2500_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1702 a_9072_4860 a_8924_5127 a_8904_4860 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1703 vccd1 a_4332_5600 a_4228_5644 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1704 vccd1 a_21740_11351 a_21652_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1705 a_37912_11045 a_32995_11784 vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X1706 a_18403_5949 a_18733_6021 a_18853_6131 vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X1707 a_33916_7864 a_35708_7864 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1708 vccd1 a_10540_11351 a_10452_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1709 vccd1 a_32236_3160 SDAC[7] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1710 vccd1 a_32565_12256 a_33284_7124 vccd1 pfet_06v0 ad=0.4005p pd=2.12u as=0.1456p ps=1.08u w=0.56u l=0.5u
X1711 a_3036_9783 a_2948_9880 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1712 vssd1 a_33500_9006 a_32964_9176 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1713 a_16926_3608 a_17004_3197 vssd1 vssd1 nfet_06v0 ad=0.1469p pd=1.085u as=0.2486p ps=2.01u w=0.565u l=0.6u
X1714 a_26513_7471 a_17640_7564 vssd1 vssd1 nfet_06v0 ad=0.2046p pd=1.81u as=0.1209p ps=0.985u w=0.465u l=0.6u
X1715 a_34818_9476 a_34678_9698 a_34054_9432 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X1716 vccd1 a_8300_11351 a_8212_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1717 a_30100_4076 a_28932_4472 a_29896_4076 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1718 vccd1 a_15940_9880 a_17696_3608 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1719 SDAC[3] a_17696_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1720 a_18044_4076 a_9632_5556 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
D83 vssd1 a_2468_4822 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1721 a_31797_8692 a_31677_9224 a_31053_9157 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1722 vssd1 a_34028_3160 a_32236_3160 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1723 a_22188_11351 a_22100_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1724 a_32040_9564 a_30240_9880 a_31100_9831 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1725 a_21871_5250 a_17640_7564 a_22289_4772 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
X1726 vccd1 a_13529_5904 a_13424_6044 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X1727 a_25248_9120 a_23599_5996 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.2344p ps=1.56u w=0.36u l=0.6u
X1728 a_26396_4032 a_26088_4076 vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X1729 SDAC[8] a_33916_7864 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1730 a_25866_11828 a_25242_11828 a_25698_11828 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1731 a_26163_11000 a_28169_10260 a_37092_7908 vssd1 nfet_06v0 ad=0.2569p pd=1.56u as=0.1312p ps=1.14u w=0.82u l=0.6u
D84 vssd1 a_2916_4822 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1732 a_10787_8312 a_10871_7864 a_10807_7909 vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X1733 vssd1 a_21392_8392 a_15324_6608 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X1734 vssd1 a_24360_9152 a_23200_4728 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X1735 vccd1 a_29132_11351 a_29044_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1736 a_17436_9831 a_17128_9880 vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
D85 XRST vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1737 a_2140_8648 a_2052_8692 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1738 vccd1 a_19916_7909 a_16569_5984 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1739 vccd1 a_13496_6366 a_2356_4118 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1740 a_3484_11784 a_3396_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1741 a_15216_7612 a_13104_7195 a_14904_7612 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X1742 a_27067_10836 a_26591_10260 vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1743 a_36609_6044 a_34420_6040 a_35737_5996 vccd1 pfet_06v0 ad=0.1079p pd=0.935u as=0.27805p ps=2.17u w=0.415u l=0.5u
X1744 vccd1 a_28040_7944 a_29263_6875 vccd1 pfet_06v0 ad=0.38705p pd=2.08u as=0.1469p ps=1.085u w=0.565u l=0.5u
X1745 a_6620_10216 a_6532_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1746 a_12197_3988 a_12077_4520 a_11453_4453 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1747 a_3720_5600 a_2468_4822 a_7156_6040 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1748 vccd1 a_4341_6296 a_4257_6744 vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1749 vssd1 a_23980_7438 a_23444_7608 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1750 vccd1 a_30163_7864 a_25784_4032 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1751 a_2356_4118 a_13496_6366 vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1752 vssd1 a_24115_5557 a_26804_7953 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1753 vccd1 a_16325_7125 a_16271_5557 vccd1 pfet_06v0 ad=0.3718p pd=2.57u as=0.2197p ps=1.365u w=0.845u l=0.5u
X1754 a_32405_11044 a_32285_11000 vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X1755 vssd1 a_24976_3608 SDAC[5] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1756 a_32680_6799 a_32279_6755 a_31623_6564 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1757 vccd1 a_17436_9831 a_17332_9880 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1758 vccd1 a_33916_7864 SDAC[8] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1759 a_36856_10748 a_34644_10744 a_35916_10304 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
D86 vssd1 a_2356_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1760 vccd1 a_30220_3160 a_28428_3160 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1761 a_5500_11784 a_5412_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1762 a_31453_10792 a_29244_9477 vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1763 vccd1 a_18403_5949 a_14975_4728 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1764 vccd1 a_21504_3608 SDAC[4] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1765 vccd1 a_2356_4118 a_9108_6423 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X1766 vssd1 a_29176_7909 a_25996_10747 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X1767 a_10871_7864 a_10751_7146 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X1768 a_6133_8693 a_5129_9040 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1769 a_37168_7612 a_35056_7195 a_36856_7612 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X1770 vccd1 CLK a_21392_8392 vccd1 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X1771 a_33992_7608 a_32565_12256 a_33768_7608 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1772 a_29440_6044 a_26916_6040 a_29128_6044 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1773 a_2936_7168 a_6252_7864 a_6148_7908 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1774 vssd1 a_17456_7080 a_17864_7080 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1775 a_16271_5557 a_16325_7125 a_16689_6040 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1517p ps=1.19u w=0.82u l=0.6u
X1776 COMP_CLK a_33916_11000 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1777 a_28169_10260 a_27439_10282 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X1778 a_30613_4772 a_30493_4728 vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X1779 a_27935_4728 a_28040_7944 vssd1 vssd1 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X1780 a_20096_10688 a_19916_7909 vccd1 vccd1 pfet_06v0 ad=0.2486p pd=2.01u as=0.35315p ps=1.96u w=0.565u l=0.5u
X1781 a_8616_5176 a_8064_5176 a_8412_5176 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1782 a_15568_5176 a_12580_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1783 a_5733_6340 a_2468_3254 vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1784 vssd1 a_17696_3608 SDAC[3] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1785 a_15881_4336 a_15464_4476 a_16257_4476 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X1786 a_15483_8723 a_15553_5512 a_15687_9176 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1722p ps=1.24u w=0.82u l=0.6u
X1787 a_5505_4476 a_1908_4118 vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X1788 a_33319_11828 a_32863_11828 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1789 a_31144_4476 a_29344_4059 a_30204_4032 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1790 vccd1 a_6496_3988 a_1908_4118 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4392p ps=1.94u w=1.22u l=0.5u
X1791 a_34104_5118 a_33511_5187 a_34840_4860 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1792 a_9196_11351 a_9108_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1793 vccd1 a_29580_11351 a_29492_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1794 a_34778_10052 a_34678_9698 a_34054_9432 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1795 a_28008_9180 a_25796_9176 a_27068_8736 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X1796 a_13994_8484 a_13370_7908 a_13846_7908 vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1797 vccd1 a_18380_11351 a_18292_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1798 a_13452_11351 a_13364_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1799 a_8412_5176 a_3696_3608 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1800 a_21180_4416 a_27776_7124 vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1801 vccd1 a_23855_11620 a_24311_11598 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1802 a_4964_3608 a_4516_3249 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X1803 vssd1 a_33916_7864 SDAC[8] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1804 a_22364_4032 a_22056_4076 vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X1805 a_26292_4076 a_25124_4472 a_26088_4076 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1806 a_10176_4860 a_8064_5176 a_9864_4860 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X1807 a_15324_6608 a_21392_8392 vssd1 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X1808 a_26507_11044 a_26031_11044 vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1809 a_31237_4772 a_31117_4728 a_30493_4728 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X1810 a_4965_4728 a_4145_3608 vccd1 vccd1 pfet_06v0 ad=0.4248p pd=1.94u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1811 a_26342_12404 a_25866_11828 a_26070_11828 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
D87 a_1908_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1812 a_33185_4472 a_30981_5996 vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1813 vssd1 a_26356_10260 a_34980_3249 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1814 a_22300_10216 a_22212_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1815 a_21252_8780 a_20084_9176 a_21048_8780 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
D88 a_3364_4822 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1816 vssd1 a_18793_9520 a_18688_9564 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X1817 a_12197_4564 a_12077_4520 a_11453_4453 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X1818 a_13860_7212 a_12692_7608 a_13656_7212 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1819 vssd1 a_13994_8484 a_14470_7908 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1820 SDAC[5] a_24976_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1821 a_6679_5176 a_6133_8693 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1822 vssd1 a_2356_4118 a_9108_6423 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1823 a_26633_7124 a_26513_7471 vccd1 vccd1 pfet_06v0 ad=0.1469p pd=1.085u as=0.38705p ps=2.08u w=0.565u l=0.5u
X1824 vccd1 a_11612_8736 a_11508_8780 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1825 vssd1 a_21504_3608 SDAC[4] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1826 a_27328_5627 a_26916_6040 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1827 vccd1 a_17416_6016 a_9532_5512 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1828 a_6496_3988 a_4964_3608 vssd1 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1829 vssd1 a_13900_4728 a_13364_4772 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1830 a_32909_11000 a_24607_5996 vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1831 a_35220_4076 a_34144_9238 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
D89 a_2468_3254 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1832 vccd1 a_15324_6608 a_27776_7124 vccd1 pfet_06v0 ad=0.2132p pd=1.34u as=0.2952p ps=1.54u w=0.82u l=0.5u
X1833 a_5584_6044 a_3060_6040 a_5272_6044 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1834 a_27215_10260 a_26591_10260 a_27067_10836 vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1835 a_3484_9783 a_3396_9880 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1836 a_3772_8736 a_3464_8780 vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X1837 a_28320_9180 a_26208_8763 a_28008_9180 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X1838 vssd1 a_28040_7944 a_27935_4728 vssd1 nfet_06v0 ad=0.1469p pd=1.085u as=0.1469p ps=1.085u w=0.565u l=0.6u
X1839 a_35608_7212 a_35056_7195 a_35404_7212 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1840 vccd1 a_20732_11784 a_20644_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1841 vssd1 a_33916_11000 COMP_CLK vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1842 a_2356_4118 a_13496_6366 vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1892p ps=1.74u w=0.43u l=0.6u
X1843 vccd1 a_13112_6044 a_13529_5904 vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X1844 a_36081_4476 a_35424_4076 vssd1 vssd1 nfet_06v0 ad=86.399994f pd=0.84u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1845 vssd1 a_21392_8392 a_15324_6608 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X1846 vccd1 a_1692_5079 a_1604_5176 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1847 a_29512_4773 a_29772_4773 vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X1848 a_26579_9432 a_26909_9432 a_27029_10030 vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1849 a_28364_7988 a_26456_8736 a_28160_7988 vssd1 nfet_06v0 ad=60.8f pd=0.7u as=79.799995f ps=0.8u w=0.38u l=0.6u
X1850 vssd1 a_37912_4773 a_37196_11045 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X1851 a_35056_7195 a_34644_7608 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X1852 a_11279_7864 a_12969_9040 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1853 vssd1 a_22157_7656 a_22277_7700 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1854 a_20496_8763 a_20084_9176 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
D90 a_2468_4822 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1855 a_29604_9880 a_29156_9521 vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X1856 a_25312_5556 a_5972_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1857 a_12244_5176 a_11796_4817 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X1858 a_24809_11448 a_24079_11044 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X1859 a_19656_7909 a_19916_7909 vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X1860 a_23072_6744 a_22660_6423 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X1861 vccd1 a_11320_6428 a_11737_6384 vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X1862 a_35220_5644 a_35100_5996 vccd1 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.22725p ps=1.91u w=0.505u l=0.5u
X1863 a_7938_7124 a_7254_7124 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1656p ps=1.28u w=0.36u l=0.5u
X1864 vssd1 a_7315_3160 a_4229_3160 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1865 vccd1 a_21504_3608 SDAC[4] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1866 a_18793_9520 a_18376_9564 a_19169_9564 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X1867 vssd1 a_19797_9477 a_20196_8000 vssd1 nfet_06v0 ad=0.2344p pd=1.56u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1868 vccd1 a_31275_6296 a_24607_5996 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1869 a_14904_7612 a_13104_7195 a_13964_7168 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1870 a_26902_12404 a_26070_11828 a_26754_11828 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1871 a_26579_9432 a_26909_9432 a_27029_9476 vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X1872 a_23855_11620 a_23231_11044 a_23707_11044 vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1873 vccd1 CLK a_21392_8392 vccd1 pfet_06v0 ad=0.428p pd=2.02u as=0.2542p ps=1.44u w=0.82u l=0.5u
X1874 a_27552_5176 a_27452_4796 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1875 vssd1 a_1908_4118 a_4480_6044 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1876 vssd1 a_33916_11000 COMP_CLK vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1877 a_35737_4428 a_22560_4292 a_36081_4476 vssd1 nfet_06v0 ad=0.1989p pd=1.465u as=86.399994f ps=0.84u w=0.36u l=0.6u
X1878 a_19656_9176 a_19052_8648 a_19432_9176 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1879 a_6496_3988 a_4964_3608 vccd1 vccd1 pfet_06v0 ad=0.2952p pd=1.54u as=0.2132p ps=1.34u w=0.82u l=0.5u
X1880 a_10752_8763 a_10340_9176 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X1881 a_22919_5557 a_23599_5996 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1882 vccd1 a_7740_11784 a_7652_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1883 a_27653_9476 a_27533_9432 a_26909_9432 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X1884 a_19808_4476 a_17284_4472 a_19496_4476 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1885 vssd1 a_21180_4416 a_29828_9559 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1886 a_7315_3160 a_7645_3160 a_7765_3758 vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1887 vssd1 a_13496_6366 a_2356_4118 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X1888 vccd1 a_33916_11000 COMP_CLK vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1889 a_32380_5870 a_28119_4728 vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1890 a_26964_8780 a_25796_9176 a_26760_8780 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1891 a_2140_10216 a_2052_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1892 a_3920_9180 a_3772_8736 a_3752_9180 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1893 SDAC[3] a_17696_3608 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1894 vssd1 a_37904_7864 a_28428_7944 vssd1 nfet_06v0 ad=0.2344p pd=1.56u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1895 a_33029_11620 a_32909_11000 a_32285_11000 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1896 vssd1 a_11279_7864 a_15492_9521 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1897 a_27676_5644 a_27236_6340 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1898 vssd1 a_21404_3160 a_21504_3608 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1899 vccd1 a_18556_4032 a_18452_4076 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1900 a_8904_4860 a_8064_5176 a_8616_5176 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1901 a_30199_6744 a_30879_6296 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1902 vssd1 a_33916_7864 SDAC[8] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1903 a_18853_6131 a_18733_6021 vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X1904 a_37092_6744 a_32481_11846 vccd1 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X1905 vccd1 a_17372_11784 a_17284_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1906 a_16140_11351 a_16052_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1907 vssd1 a_22560_4292 a_31248_9564 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1908 a_2936_7168 a_4257_6744 vccd1 vccd1 pfet_06v0 ad=0.4248p pd=1.94u as=0.4972p ps=3.14u w=1.13u l=0.5u
X1909 vccd1 a_24092_10216 a_24004_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1910 vccd1 a_22157_7656 a_22277_7124 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X1911 a_15324_6608 a_21392_8392 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1912 a_26163_11000 a_36972_7864 a_36884_8312 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
D91 COMP_OUT vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
D92 a_2356_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1913 a_34678_9698 a_35090_9432 a_35210_9476 vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1914 a_24976_3608 a_24876_3160 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1915 a_25629_4728 a_23652_7608 vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1916 a_27691_10835 a_27215_10260 a_27439_10282 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X1917 vccd1 a_4828_10216 a_4740_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1918 vccd1 a_21180_4416 a_21092_4472 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X1919 vssd1 a_8086_7700 a_8562_7699 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X1920 vccd1 a_35336_4816 a_35232_4860 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1921 vssd1 a_21180_4416 a_22660_6423 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X1922 vccd1 a_37513_5984 a_36833_6044 vccd1 pfet_06v0 ad=0.3276p pd=1.62u as=0.2028p ps=1.3u w=0.78u l=0.5u
X1923 a_7168_8312 a_6756_7991 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X1924 a_10100_5556 a_9980_5870 vccd1 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X1925 vssd1 a_4573_4728 a_4693_4772 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1926 vssd1 a_1908_4118 a_10528_6428 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1927 SDAC[8] a_33916_7864 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1928 vssd1 a_22560_4292 a_32995_4852 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=0.134p ps=1.1u w=0.36u l=0.6u
X1929 a_2140_9783 a_2052_9880 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1930 a_35834_10052 a_35714_9432 a_35090_9432 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1931 a_35834_9476 a_35714_9432 a_35090_9432 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X1932 SDAC[4] a_21504_3608 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1933 a_12864_9180 a_10340_9176 a_12552_9180 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1934 vccd1 a_9717_4416 a_9633_4006 vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X1935 a_22919_5557 a_17640_7564 a_23107_5557 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1936 a_33407_5231 a_32507_4728 vccd1 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.29465p ps=1.74u w=0.505u l=0.5u
X1937 a_12244_5176 a_11796_4817 vssd1 vssd1 nfet_06v0 ad=0.2178p pd=1.87u as=0.153p ps=1.195u w=0.495u l=0.6u
X1938 a_27111_11598 a_26655_11620 a_26879_11044 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X1939 vccd1 a_19972_9476 a_16365_5984 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1940 vccd1 a_17864_7080 a_17368_7124 vccd1 pfet_06v0 ad=0.4005p pd=2.12u as=0.3172p ps=1.74u w=1.22u l=0.5u
X1941 vssd1 a_28428_7944 a_36084_6377 vssd1 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
D93 a_1908_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1942 vccd1 a_35708_11000 a_33916_11000 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1943 vssd1 a_17696_3608 SDAC[3] vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1944 a_3932_11351 a_3844_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X1945 vssd1 a_12600_7909 a_9980_5870 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X1946 vccd1 a_2356_4118 a_2500_4472 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X1947 vccd1 a_33094_5892 a_2468_3254 vccd1 pfet_06v0 ad=0.4941p pd=2.03u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1948 vccd1 a_23420_11784 a_23332_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1949 a_33132_6744 a_32680_6799 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.45p ps=2.02u w=0.78u l=0.5u
X1950 a_30199_6744 a_30471_6296 a_30387_6744 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X1951 vssd1 a_32995_11784 a_32863_11828 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X1952 vccd1 a_36856_10748 a_37273_10608 vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X1953 SDAC[6] a_28428_3160 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1954 vssd1 a_19916_7909 a_16569_5984 vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1955 a_10072_6744 a_9108_6423 a_9868_6744 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
D94 vssd1 a_2356_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1956 a_29545_5904 a_29128_6044 a_29921_6044 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X1957 a_26302_11828 a_25866_11828 a_26070_11828 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X1958 a_3820_5644 a_3720_5600 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X1959 a_19913_4336 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X1960 a_34888_9152 a_32565_12256 vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
D95 a_1908_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X1961 a_23295_10052 a_22671_9476 a_23147_9476 vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1962 a_12992_3988 a_12892_3944 vssd1 vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X1963 a_11860_7908 a_12188_7864 a_9768_6574 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1964 a_29128_6044 a_26916_6040 a_28188_5600 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X1965 a_12220_3205 a_15881_4336 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X1966 a_33916_7864 a_35708_7864 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1967 a_31465_5512 a_32404_7864 vccd1 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X1968 a_8157_6296 a_5909_7125 vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X1969 a_17114_3608 a_17004_3197 a_16926_3608 vccd1 pfet_06v0 ad=0.4087p pd=1.89u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1970 a_24976_3608 a_24876_3160 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1971 a_31509_7864 a_22848_5176 a_31844_6040 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X1972 a_21203_5949 a_21533_6021 a_21653_6131 vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
D96 vssd1 a_3364_4822 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X1973 a_32964_9176 a_28040_7944 a_30488_9710 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1974 a_34144_9238 a_30913_5557 vssd1 vssd1 nfet_06v0 ad=0.2569p pd=1.56u as=0.2244p ps=1.9u w=0.51u l=0.6u
X1975 a_4712_4476 a_2912_4059 a_3772_4032 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X1976 vccd1 a_1692_11351 a_1604_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X1977 vccd1 a_23980_7438 a_23652_7608 vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.4248p ps=1.94u w=1.13u l=0.5u
X1978 a_22560_4292 a_25312_5556 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X1979 a_23771_9476 a_23295_10052 a_23519_9476 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X1980 a_11612_8736 a_11304_8780 vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X1981 a_3036_7212 a_2936_7168 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X1982 a_5129_9040 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X1983 vccd1 a_18536_10720 a_15383_8679 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X1984 a_12220_3205 a_15881_4336 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1985 a_22364_4032 a_22056_4076 vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X1986 a_6887_4773 a_3364_4822 vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X1987 vssd1 a_1908_4118 a_11760_9180 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X1988 SDAC[7] a_32236_3160 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1989 a_24543_6040 a_21871_6818 a_24115_5557 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X1990 vccd1 a_4488_7612 a_4905_7472 vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X1991 a_11864_5644 a_10900_6040 a_11660_5644 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X1992 vccd1 a_29244_9477 a_29156_9521 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1993 vssd1 a_28040_7944 a_32932_7908 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1148p ps=1.1u w=0.82u l=0.6u
X1994 vccd1 a_2356_4118 a_17284_4472 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X1995 a_16364_6296 a_16694_6296 a_16814_6340 vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X1996 a_15324_6608 a_21392_8392 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1997 a_37912_4773 a_33768_7608 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X1998 a_17696_3608 a_15940_9880 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X1999 vssd1 a_12220_3205 a_12132_3249 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2000 vccd1 a_15483_8723 a_19089_6744 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2001 a_4277_6340 a_2468_3254 vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2002 a_31623_6564 a_32279_6755 a_32175_6799 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.1313p ps=1.025u w=0.505u l=0.5u
X2003 a_23868_11784 a_23780_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2004 a_33916_11000 a_35708_11000 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2005 a_3720_5600 a_5713_6744 vccd1 vccd1 pfet_06v0 ad=0.4248p pd=1.94u as=0.4972p ps=3.14u w=1.13u l=0.5u
D97 vssd1 COMP_OUT diode_nd2ps_06v0 pj=1.86u area=0.2052p
D98 a_1908_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2006 a_27533_9432 a_26293_6341 vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X2007 a_22296_9180 a_20496_8763 a_21356_8736 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2008 vssd1 a_30163_7864 a_25784_4032 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2009 a_15030_7908 a_14198_8402 a_14862_7908 vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2010 a_34840_4860 a_33912_5231 a_34672_4860 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2011 a_29440_6044 a_27328_5627 a_29128_6044 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X2012 vssd1 a_33916_7864 SDAC[8] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2013 a_13653_10260 a_13533_10792 a_12909_10725 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2014 a_30996_9880 a_22560_4292 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X2015 vssd1 a_20495_6296 a_20028_7080 vssd1 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2016 vssd1 a_7203_6296 a_4341_6296 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2017 a_28428_3160 a_30220_3160 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2018 a_15324_6608 a_21392_8392 vssd1 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X2019 a_32977_3989 a_29739_6744 vccd1 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2020 vccd1 a_2916_4822 a_25159_7125 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
D99 vssd1 a_3364_4822 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2021 SDAC[2] a_15568_5176 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2022 vccd1 a_21203_5949 a_20127_4728 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2023 a_7516_8312 a_7416_8142 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X2024 vccd1 a_31144_4476 a_31561_4336 vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X2025 a_10988_11351 a_10900_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2026 a_21392_8392 CLK vccd1 vccd1 pfet_06v0 ad=0.2542p pd=1.44u as=0.2542p ps=1.44u w=0.82u l=0.5u
X2027 a_18044_4076 a_9632_5556 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2028 a_28336_6044 a_28188_5600 a_28168_6044 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2029 a_5272_6044 a_3060_6040 a_4332_5600 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X2030 a_32384_6384 a_21180_4416 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
D100 vssd1 a_2468_3254 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2031 a_32872_6686 a_32279_6755 a_33608_6428 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2032 a_13664_4059 a_13252_4472 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2033 a_8748_11351 a_8660_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2034 a_7203_6296 a_7533_6296 a_7653_6894 vccd1 pfet_06v0 ad=0.3456p pd=2.64u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2035 a_26902_12404 a_26070_11828 a_26734_12404 vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2036 vssd1 a_1908_4118 a_14672_4476 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2037 SDAC[5] a_24976_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2038 vccd1 a_24876_3160 a_24976_3608 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2039 vccd1 a_17932_11351 a_17844_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2040 vssd1 a_29604_9880 a_32964_10791 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2041 a_29772_4773 a_29739_6744 a_33185_4472 vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2042 a_6036_4772 a_4145_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2043 a_37649_10748 a_22560_4292 vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X2044 a_19432_8692 a_18760_8692 vccd1 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4005p ps=2.12u w=1.22u l=0.5u
X2045 a_33029_11044 a_32909_11000 a_32285_11000 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X2046 SDAC[4] a_21504_3608 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2047 vssd1 a_25312_5556 a_22560_4292 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2048 a_10527_7124 a_9903_7124 a_10359_7124 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2049 vssd1 a_34888_9152 a_32404_7864 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X2050 vccd1 a_30668_7577 a_31226_7124 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2051 a_20523_7608 a_20403_7098 a_18828_9199 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2052 a_22085_4772 a_20495_6296 a_21891_4772 vssd1 nfet_06v0 ad=0.1722p pd=1.24u as=0.1517p ps=1.19u w=0.82u l=0.6u
X2053 a_21871_5250 a_19052_8648 vccd1 vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X2054 vccd1 a_7516_10216 a_7428_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2055 a_22277_7700 a_22157_7656 a_21533_7589 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X2056 a_17864_7080 a_17640_7564 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.218p ps=1.52u w=0.36u l=0.6u
X2057 vssd1 a_31955_11000 a_30879_6296 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2058 a_29344_4059 a_28932_4472 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2059 a_32395_10744 a_28428_7944 a_30668_7577 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2060 vssd1 a_17864_8648 a_16824_9710 vssd1 nfet_06v0 ad=0.218p pd=1.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2061 a_5584_6044 a_3472_5627 a_5272_6044 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X2062 a_5909_7125 a_4905_7472 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2063 SDAC[6] a_28428_3160 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2064 vccd1 a_4828_11784 a_4740_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2065 a_28084_5644 a_26916_6040 a_27880_5644 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2066 vssd1 a_21392_8392 a_15324_6608 vssd1 nfet_06v0 ad=0.1261p pd=1.005u as=0.1261p ps=1.005u w=0.485u l=0.6u
X2067 SDAC[4] a_21504_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2068 vccd1 a_24249_9880 a_35336_4816 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2069 a_13364_4772 a_2468_4822 a_11560_5600 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2070 a_27748_7864 a_28428_7944 a_28364_7988 vssd1 nfet_06v0 ad=0.1672p pd=1.64u as=60.8f ps=0.7u w=0.38u l=0.6u
X2071 a_30668_7577 a_28428_7944 vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X2072 a_18688_9564 a_16164_9559 a_18376_9564 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2073 vssd1 a_1908_4118 a_14112_7612 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2074 a_5024_9180 a_2912_8763 a_4712_9180 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X2075 a_18556_4032 a_18248_4076 vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
D101 vssd1 a_1908_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2076 vccd1 a_26655_11620 a_27111_11598 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2077 a_28008_9180 a_26208_8763 a_27068_8736 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2078 a_7765_3758 a_7645_3160 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X2079 vssd1 a_24976_3608 SDAC[5] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2080 vccd1 a_7964_10216 a_7876_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2081 a_9717_4416 a_15254_7908 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X2082 a_3752_9180 a_2912_8763 a_3464_8780 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2083 vccd1 a_4905_7472 a_4800_7612 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X2084 vccd1 a_4380_11351 a_4292_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2085 a_18556_4032 a_18248_4076 vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X2086 a_27378_12403 a_26902_12404 a_27126_11850 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X2087 vccd1 a_11279_7864 a_16625_8312 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2088 a_29921_6044 a_22560_4292 vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X2089 vssd1 a_21180_4416 a_26916_6040 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2090 vccd1 a_2468_3254 a_23980_7438 vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X2091 a_2688_7195 a_2276_7608 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
D102 vssd1 a_1908_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2092 vccd1 a_29176_7909 a_25996_10747 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2093 vssd1 a_24809_11448 a_34292_8648 vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X2094 a_5972_3608 a_5524_3249 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X2095 vssd1 a_25374_11784 a_25242_11828 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X2096 vccd1 a_26456_8736 a_27748_7864 vccd1 pfet_06v0 ad=0.1391p pd=1.055u as=0.1391p ps=1.055u w=0.535u l=0.5u
X2097 SDAC[3] a_17696_3608 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2098 vccd1 a_3228_3228 a_3140_3272 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2099 a_22277_7124 a_22157_7656 a_21533_7589 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2100 vccd1 a_7484_5512 a_7380_5556 vccd1 pfet_06v0 ad=0.5978p pd=3.42u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2101 a_16715_7608 a_14567_4728 a_13900_4728 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2102 a_15483_8723 a_15553_5512 vccd1 vccd1 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2103 vccd1 a_22188_11351 a_22100_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2104 a_12172_5600 a_11864_5644 vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X2105 vccd1 a_27753_4336 a_27648_4476 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X2106 a_8562_7699 a_8086_7700 a_8310_7146 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.3705p ps=2.77u w=0.365u l=0.6u
X2107 a_33172_8692 a_30668_7577 vccd1 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.5978p ps=3.42u w=1.22u l=0.5u
X2108 a_31677_9224 a_22932_4728 vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X2109 a_36972_7864 a_37780_9568 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2344p ps=1.56u w=0.82u l=0.6u
X2110 a_15356_11784 a_15268_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2111 vssd1 a_35336_4816 a_35232_4860 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2112 a_4693_4772 a_4573_4728 a_3949_4728 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.369p ps=2.77u w=0.36u l=0.6u
X2113 a_8064_5176 a_7652_4855 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2114 a_31955_11000 a_32285_11000 a_32405_11044 vssd1 nfet_06v0 ad=0.3705p pd=2.77u as=43.8f ps=0.605u w=0.365u l=0.6u
X2115 a_34832_4059 a_34420_4472 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2116 vccd1 a_28428_3160 SDAC[6] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2117 a_4069_5326 a_3949_4728 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X2118 vssd1 a_21180_4416 a_34420_6040 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
D103 a_2468_3254 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2119 vssd1 a_27753_4336 a_27648_4476 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
D104 a_1908_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2120 a_12552_9180 a_10340_9176 a_11612_8736 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X2121 vccd1 a_22713_9040 a_22608_9180 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X2122 vccd1 a_34104_6384 a_34000_6428 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2123 a_20609_5176 a_19524_11448 vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X2124 a_13424_6044 a_10900_6040 a_13112_6044 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2125 a_8007_6040 a_3364_4822 vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2126 a_4165_3204 a_2468_3254 vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2127 a_11612_8736 a_11304_8780 vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X2128 vccd1 a_15324_6608 a_27776_7124 vccd1 pfet_06v0 ad=0.367p pd=1.92u as=0.2952p ps=1.54u w=0.82u l=0.5u
X2129 a_18948_8692 a_18828_9199 a_18760_8692 vccd1 pfet_06v0 ad=0.1456p pd=1.08u as=0.2464p ps=2u w=0.56u l=0.5u
X2130 vccd1 a_24976_3608 SDAC[5] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2131 vccd1 a_23932_6695 a_23828_6744 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2132 vccd1 a_8086_7700 a_8542_7146 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2133 a_36833_4476 a_34832_4059 a_36609_4476 vccd1 pfet_06v0 ad=0.1826p pd=1.71u as=0.1079p ps=0.935u w=0.415u l=0.5u
X2134 a_2588_6647 a_2500_6744 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2135 vccd1 a_28040_7944 a_31465_5512 vccd1 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2136 vccd1 a_16924_11784 a_16836_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2137 a_3668_8780 a_2500_9176 a_3464_8780 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2138 a_27236_6340 a_27116_6296 a_27028_6340 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2139 a_7068_10216 a_6980_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2140 SDAC[5] a_24976_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2141 vccd1 a_23644_10216 a_23556_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2142 a_6065_6044 a_1908_4118 vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X2143 vssd1 a_2356_4118 a_3060_6040 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2144 a_31573_10260 a_31453_10792 a_30829_10725 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2145 a_11324_10216 a_11236_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2146 a_37912_3205 a_22932_4728 vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X2147 vccd1 a_12556_4773 a_12468_4817 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
D105 a_2356_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2148 a_27609_11448 a_26879_11044 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X2149 a_17456_7080 a_18940_7080 vccd1 vccd1 pfet_06v0 ad=0.4334p pd=2.85u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2150 vccd1 a_3548_7168 a_3444_7212 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2151 vccd1 a_25629_4728 a_25749_5348 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2152 vccd1 a_34678_9698 a_34778_10052 vccd1 pfet_06v0 ad=0.1656p pd=1.28u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2153 a_19432_9176 a_18760_8692 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X2154 a_26208_8763 a_25796_9176 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2155 vccd1 a_32236_3160 SDAC[7] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2156 a_10204_11784 a_10116_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D106 a_2916_4822 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2157 a_21653_6131 a_21533_6021 vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X2158 vssd1 a_30668_7577 a_27935_4728 vssd1 nfet_06v0 ad=0.2486p pd=2.01u as=0.1469p ps=1.085u w=0.565u l=0.6u
X2159 a_32405_11598 a_32285_11000 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X2160 a_5713_6744 a_2468_3254 vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X2161 a_12864_9180 a_10752_8763 a_12552_9180 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X2162 a_1692_5512 a_1604_5556 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2163 vccd1 a_21392_8392 a_15324_6608 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2164 a_19524_11448 a_19076_11089 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X2165 a_26655_11620 a_26031_11044 a_26507_11044 vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2166 vccd1 a_17696_3608 SDAC[3] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2167 a_25775_7608 a_2916_4822 a_23052_7564 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X2168 vccd1 a_9196_11351 a_9108_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2169 vccd1 a_28428_3160 SDAC[6] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2170 a_9864_4860 a_8064_5176 a_8924_5127 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2171 a_30924_11351 a_30836_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2172 a_27564_6296 a_30471_6296 vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X2173 a_9768_6574 a_9633_4006 vccd1 vccd1 pfet_06v0 ad=0.4248p pd=1.94u as=0.4972p ps=3.14u w=1.13u l=0.5u
X2174 a_14295_5176 a_14975_4728 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2175 a_8616_5176 a_7652_4855 a_8412_5176 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2176 vccd1 a_13452_11351 a_13364_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2177 vssd1 a_27776_7124 a_21180_4416 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2178 SDAC[8] a_33916_7864 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2179 a_5689_5904 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X2180 a_21871_6818 a_17004_3197 vccd1 vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X2181 vssd1 a_21392_8392 a_15324_6608 vssd1 nfet_06v0 ad=0.2134p pd=1.85u as=0.1261p ps=1.005u w=0.485u l=0.6u
X2182 a_17820_11784 a_17732_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D107 a_2356_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2183 a_35428_3608 a_34980_3249 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X2184 a_10276_6744 a_9108_6423 a_10072_6744 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2185 vccd1 a_3036_10216 a_2948_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2186 a_16814_6340 a_16694_6296 vssd1 vssd1 nfet_06v0 ad=43.8f pd=0.605u as=0.282625p ps=1.87u w=0.365u l=0.6u
X2187 vccd1 a_13496_6366 a_2356_4118 vccd1 pfet_06v0 ad=0.367p pd=1.92u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2188 vssd1 a_20127_4728 a_20063_4773 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2189 vssd1 a_24876_3160 a_24976_3608 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2190 vccd1 a_37196_11045 a_36884_8312 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.44955p ps=1.955u w=1.215u l=0.5u
X2191 vccd1 a_8028_8263 a_7924_8312 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2192 a_3260_8780 a_3140_3272 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X2193 a_15503_9176 a_15383_8679 vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2194 a_35056_10331 a_34644_10744 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2195 a_23927_5557 a_24607_5996 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
D108 a_2356_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2196 a_14862_7908 a_14198_8402 vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2197 a_30100_4076 a_22560_4292 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X2198 a_34672_4860 a_22560_4292 vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.2016p ps=1.48u w=0.36u l=0.6u
X2199 a_12113_6428 a_1908_4118 vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X2200 SDAC[5] a_24976_3608 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2201 vssd1 a_24976_3608 SDAC[5] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2202 vccd1 a_28348_11784 a_28260_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2203 vccd1 a_4712_4476 a_5129_4336 vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X2204 vccd1 a_37196_11045 a_37108_11089 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X2205 a_17368_8692 a_16365_5984 a_16824_9710 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.3172p ps=1.74u w=1.22u l=0.5u
X2206 a_3240_7212 a_2688_7195 a_3036_7212 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2207 vccd1 a_21504_3608 SDAC[4] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2208 a_16924_9880 a_16824_9710 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2209 a_6396_11784 a_6308_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2210 vccd1 a_33916_11000 COMP_CLK vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2211 a_9532_10216 a_9444_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2212 a_2140_11351 a_2052_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2213 a_16365_5984 a_19972_9476 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.4941p ps=2.03u w=1.22u l=0.5u
X2214 a_2912_8763 a_2500_9176 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2215 a_10652_11784 a_10564_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2216 a_30725_5557 a_30981_5996 a_30913_5557 vccd1 pfet_06v0 ad=0.37665p pd=1.835u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2217 a_28168_6044 a_27328_5627 a_27880_5644 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2218 vssd1 a_24607_5996 a_24543_6040 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2219 a_35424_4076 a_34832_4059 a_35220_4076 vccd1 pfet_06v0 ad=0.19315p pd=1.27u as=0.1313p ps=1.025u w=0.505u l=0.5u
X2220 a_33608_6428 a_32680_6799 a_33440_6428 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2221 a_14616_9477 a_14876_9477 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X2222 vccd1 a_27748_7864 a_17456_8648 vccd1 pfet_06v0 ad=0.4268p pd=2.175u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2223 a_7653_6894 a_7533_6296 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X2224 a_14672_4476 a_14524_4032 a_14504_4476 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2225 a_2468_3254 a_33094_5892 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2226 vccd1 a_16926_3608 a_20420_6087 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X2227 vccd1 a_5972_3608 a_25312_5556 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2228 SDAC[2] a_15568_5176 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2229 vccd1 a_4828_9783 a_4740_9880 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2230 vccd1 a_22296_9180 a_22713_9040 vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X2231 a_10359_7124 a_9903_7124 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.1116p ps=0.98u w=0.36u l=0.5u
X2232 a_19496_4476 a_17284_4472 a_18556_4032 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X2233 vccd1 a_14904_7612 a_15321_7472 vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X2234 a_21392_8392 CLK vccd1 vccd1 pfet_06v0 ad=0.2542p pd=1.44u as=0.3608p ps=2.52u w=0.82u l=0.5u
X2235 vssd1 a_2356_4118 a_10900_6040 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2236 a_33916_11000 a_35708_11000 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2237 a_27856_11828 a_27126_11850 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
D109 vssd1 a_2356_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2238 vccd1 a_3484_10216 a_3396_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2239 vccd1 a_8157_6296 a_8277_6916 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2240 vssd1 a_31117_4728 a_31237_4772 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2241 a_24115_5557 a_17640_7564 a_24135_6040 vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2242 a_30488_9710 a_30668_7577 a_32964_9176 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2243 a_14540_8648 a_11285_4773 vssd1 vssd1 nfet_06v0 ad=0.2569p pd=1.56u as=0.2244p ps=1.9u w=0.51u l=0.6u
X2244 a_31304_3205 a_24607_5996 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X2245 vccd1 a_35916_10304 a_35812_10348 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2246 a_24809_11448 a_24079_11044 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X2247 a_32855_4996 a_33616_4816 a_33407_5231 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=94.5f ps=0.885u w=0.36u l=0.6u
X2248 a_23196_10216 a_23108_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2249 vssd1 a_2356_4118 a_6756_7991 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2250 vssd1 a_27564_6296 a_27028_6340 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2251 vccd1 a_23363_11000 a_23231_11044 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2252 a_9980_10216 a_9892_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D110 vssd1 a_2468_3254 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2253 vssd1 a_10428_5870 a_9892_6040 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2254 vccd1 a_7050_7124 a_7486_7124 vccd1 pfet_06v0 ad=0.1656p pd=1.28u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2255 a_4604_8215 a_4516_8312 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2256 a_13529_5904 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X2257 vccd1 a_19612_11784 a_19524_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2258 a_30204_4032 a_29896_4076 vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X2259 a_22076_11784 a_21988_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2260 a_35608_10348 a_35056_10331 a_35404_10348 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2261 vssd1 a_22713_9040 a_22608_9180 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X2262 a_17904_8312 a_18236_7864 a_14540_8648 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2263 a_20495_6296 a_20196_8000 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.35315p ps=1.96u w=1.22u l=0.5u
D111 a_2468_3254 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2264 vccd1 a_30252_11784 a_30164_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2265 vccd1 a_21392_8392 a_15324_6608 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2266 a_6260_5176 a_6140_4728 a_4965_4728 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4248p ps=1.94u w=1.22u l=0.5u
X2267 a_19808_4476 a_17696_4059 a_19496_4476 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X2268 a_16625_8312 a_15383_8679 a_12860_7909 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.3159p ps=1.735u w=1.215u l=0.5u
D112 vssd1 a_2356_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2269 a_4380_9783 a_4292_9880 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2270 vssd1 a_32384_6384 a_32279_6755 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2271 a_19361_6296 a_19913_4336 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2272 a_2356_4118 a_13496_6366 vssd1 vssd1 nfet_06v0 ad=0.1118p pd=0.95u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2273 vccd1 a_30220_3160 a_28428_3160 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2274 a_21252_8780 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X2275 a_34104_6384 a_30387_6744 vssd1 vssd1 nfet_06v0 ad=0.2112p pd=1.84u as=0.2112p ps=1.84u w=0.48u l=0.6u
X2276 a_37092_9476 a_36084_6377 vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2277 vccd1 a_12600_7909 a_9980_5870 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2278 a_5909_7125 a_4905_7472 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2279 a_23721_4336 a_23304_4476 a_24097_4476 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X2280 vccd1 a_21404_3160 a_21504_3608 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2281 a_22560_4292 a_25312_5556 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2282 a_12969_9040 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X2283 vssd1 a_1908_4118 a_27216_9180 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2284 a_21852_4076 a_21752_4032 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X2285 vccd1 a_8188_11784 a_8100_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2286 a_15464_4476 a_13252_4472 a_14524_4032 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X2287 a_15568_5176 a_12580_3608 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2288 a_29804_10216 a_29716_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2289 a_7068_9783 a_6980_9880 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2290 a_18172_7908 a_16325_7125 a_14540_8648 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.2569p ps=1.56u w=0.82u l=0.6u
X2291 vccd1 a_12444_11784 a_12356_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2292 vssd1 a_2356_4118 a_13252_4472 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2293 vccd1 a_16140_11351 a_16052_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2294 a_30204_4032 a_29896_4076 vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X2295 a_31275_6296 a_31623_6564 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.44p ps=2.88u w=1u l=0.5u
X2296 a_1692_11784 a_1604_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
D113 a_2468_4822 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2297 vccd1 a_25368_10720 a_15737_5996 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2298 vccd1 a_35714_9432 a_35834_10052 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2299 a_24976_3608 a_24876_3160 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2300 a_35668_6044 a_34832_5627 a_35424_5644 vssd1 nfet_06v0 ad=62.1f pd=0.705u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2301 a_23072_6744 a_22660_6423 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2302 a_21180_4416 a_27776_7124 vccd1 vccd1 pfet_06v0 ad=0.4392p pd=1.94u as=0.367p ps=1.92u w=1.22u l=0.5u
X2303 a_15568_5176 a_12580_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2304 vccd1 a_8968_7996 a_9385_7952 vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X2305 a_1692_7080 a_1604_7124 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2306 vssd1 a_32565_12256 a_33096_7124 vssd1 nfet_06v0 ad=0.218p pd=1.52u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2307 vccd1 a_6496_3988 a_1908_4118 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2308 SC a_35708_9001 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2309 vccd1 a_9385_7952 a_9280_7996 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X2310 vccd1 a_29512_4773 a_22803_9432 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.5368p ps=3.32u w=1.22u l=0.5u
D114 a_2468_3254 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2311 a_35714_9432 a_30549_5557 vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2312 vccd1 a_19797_9477 a_19972_9476 vccd1 pfet_06v0 ad=0.4941p pd=2.03u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2313 a_11215_7909 a_2916_4822 a_10787_8312 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X2314 vccd1 a_31465_5512 a_31341_5557 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.37665p ps=1.835u w=1.215u l=0.5u
X2315 a_13112_6044 a_10900_6040 a_12172_5600 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X2316 vssd1 a_29604_9880 a_32395_10744 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2317 vccd1 a_17696_3608 SDAC[3] vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2318 vccd1 a_3932_11351 a_3844_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2319 a_16824_9710 a_16365_5984 a_17576_9176 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2320 a_15324_6608 a_21392_8392 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
D115 a_2916_4822 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2321 a_24540_11784 a_24452_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2322 a_15776_4476 a_13664_4059 a_15464_4476 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X2323 vccd1 a_3036_11784 a_2948_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2324 a_8542_7146 a_8086_7700 a_8310_7146 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3456p ps=2.64u w=0.36u l=0.5u
X2325 a_27328_5627 a_26916_6040 vccd1 vccd1 pfet_06v0 ad=0.3806p pd=2.61u as=0.2249p ps=1.385u w=0.865u l=0.5u
X2326 a_3548_7168 a_3240_7212 vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X2327 a_6252_7864 a_16108_3228 vssd1 vssd1 nfet_06v0 ad=0.1248p pd=1u as=0.2112p ps=1.84u w=0.48u l=0.6u
X2328 vccd1 a_28428_3160 SDAC[6] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2329 vccd1 a_25312_5556 a_22560_4292 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2330 vssd1 a_13496_6366 a_2356_4118 vssd1 nfet_06v0 ad=0.1892p pd=1.74u as=0.1118p ps=0.95u w=0.43u l=0.6u
X2331 a_10360_6428 a_9520_6744 a_10072_6744 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2332 vssd1 a_2468_3254 a_16715_7608 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2333 a_8028_8263 a_7720_8312 vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X2334 a_27452_4796 a_28119_4728 a_28055_4773 vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2335 a_3548_7168 a_3240_7212 vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X2336 vccd1 a_12220_3205 a_15057_5557 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2337 a_4228_5644 a_3060_6040 a_4024_5644 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2338 a_11560_5600 a_12916_5176 a_13364_4772 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2339 a_17576_7608 a_17456_7080 vssd1 vssd1 nfet_06v0 ad=0.1312p pd=1.14u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2340 vccd1 a_34104_5118 a_33912_5231 vccd1 pfet_06v0 ad=0.2222p pd=1.89u as=0.2424p ps=1.465u w=0.505u l=0.5u
X2341 vssd1 a_35708_7864 a_33916_7864 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
D116 vssd1 a_2468_4822 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2342 vssd1 a_31275_6296 a_24607_5996 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2343 a_25749_5348 a_25629_4728 a_25005_4728 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2344 a_18536_4476 a_17696_4059 a_18248_4076 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2345 a_1692_6647 a_1604_6744 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2346 vccd1 a_6172_10216 a_6084_10260 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2347 a_35714_9432 a_30549_5557 vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X2348 vccd1 a_2356_4118 a_6756_7991 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2349 a_1692_3511 a_1604_3608 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2350 vssd1 a_34104_6384 a_34000_6428 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
D117 vssd1 a_16108_3228 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2351 a_14908_11784 a_14820_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2352 a_17640_7564 a_15553_5512 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2353 vccd1 a_22000_9432 a_21404_3160 vccd1 pfet_06v0 ad=0.35315p pd=1.96u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2354 SDAC[5] a_24976_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2355 vccd1 a_30163_4728 a_25839_7564 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2356 a_4145_3608 a_4229_3160 a_4165_3204 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2357 vccd1 a_19052_8648 a_18948_8692 vccd1 pfet_06v0 ad=0.4005p pd=2.12u as=0.1456p ps=1.08u w=0.56u l=0.5u
X2358 a_26556_8780 a_26456_8736 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2359 a_13424_6044 a_11312_5627 a_13112_6044 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
D118 vssd1 a_16108_3228 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2360 vssd1 a_12579_10653 a_11740_9500 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2361 a_17416_6016 a_17676_5512 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X2362 vssd1 a_31465_5512 a_37435_3204 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2363 vssd1 a_2356_4118 a_2276_7608 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2364 vccd1 a_24540_9783 a_24452_9880 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2365 vssd1 a_35714_9432 a_35834_9476 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2366 vssd1 a_1908_4118 a_9072_4860 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2367 vccd1 a_9864_4860 a_10281_4816 vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X2368 vccd1 a_13533_10792 a_13653_10260 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2369 vccd1 a_2916_4822 a_27847_5176 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2370 a_33487_11828 a_32863_11828 a_33339_12404 vssd1 nfet_06v0 ad=0.369p pd=2.77u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2371 vccd1 a_21392_8392 a_15324_6608 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2372 a_35056_7195 a_34644_7608 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2373 vccd1 a_3484_11784 a_3396_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
D119 a_2356_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2374 a_32995_4852 a_32855_4996 a_32507_4728 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.176p ps=1.68u w=0.4u l=0.6u
X2375 a_4257_6744 a_2468_3254 vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
X2376 a_9532_9783 a_9444_9880 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2377 a_25368_10720 a_20868_5556 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X2378 a_16271_5557 a_16569_5984 vccd1 vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X2379 a_25125_5326 a_25005_4728 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X2380 vccd1 a_8924_5127 a_8820_5176 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2381 vccd1 a_12969_9040 a_12864_9180 vccd1 pfet_06v0 ad=0.29465p pd=1.74u as=0.1313p ps=1.025u w=0.505u l=0.5u
X2382 a_27648_4476 a_25124_4472 a_27336_4476 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2383 vccd1 a_5500_11784 a_5412_11828 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2384 a_35232_4860 a_33616_4816 a_34104_5118 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2385 vssd1 a_25839_7564 a_25775_7608 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2386 vssd1 a_3619_4728 a_3160_4032 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
D120 a_3364_4822 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2387 vssd1 a_25289_6384 a_25184_6428 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X2388 SDAC[6] a_28428_3160 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2389 vssd1 a_15568_5176 SDAC[2] vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2390 vccd1 a_31465_5512 a_27564_6296 vccd1 pfet_06v0 ad=0.4972p pd=3.14u as=0.2938p ps=1.65u w=1.13u l=0.5u
X2391 vccd1 a_10988_11351 a_10900_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2392 vccd1 a_20495_6296 a_20411_6760 vccd1 pfet_06v0 ad=0.2561p pd=1.505u as=0.2561p ps=1.505u w=0.985u l=0.5u
X2393 a_12969_9040 a_12552_9180 a_13345_9180 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X2394 a_34000_6428 a_32384_6384 a_32872_6686 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2395 a_17318_6562 a_17730_6296 a_17870_6916 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2396 vccd1 a_8748_11351 a_8660_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2397 SDAC[5] a_24976_3608 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2398 a_6496_3988 a_4964_3608 vccd1 vccd1 pfet_06v0 ad=0.2952p pd=1.54u as=0.3608p ps=2.52u w=0.82u l=0.5u
X2399 a_25100_11351 a_25012_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2400 a_33593_4472 a_24809_11448 a_29772_4773 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.2119p ps=1.335u w=0.815u l=0.6u
X2401 a_14504_4476 a_13664_4059 a_14216_4076 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2402 a_4380_11784 a_4292_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2403 vccd1 a_25248_9120 a_24876_3160 vccd1 pfet_06v0 ad=0.35315p pd=1.96u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2404 a_15687_9176 a_6252_7864 a_15503_9176 vssd1 nfet_06v0 ad=0.1722p pd=1.24u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2405 a_29896_4076 a_29344_4059 a_29692_4076 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2406 vccd1 a_26579_9432 a_24435_7098 vccd1 pfet_06v0 ad=0.379p pd=2.37u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2407 vssd1 a_11285_4773 a_11796_4817 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2408 a_11737_6384 a_11320_6428 a_12113_6428 vssd1 nfet_06v0 ad=0.176p pd=1.68u as=0.134p ps=1.1u w=0.4u l=0.6u
X2409 a_10035_7080 a_9385_7952 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2410 a_18354_6296 a_14533_5557 vccd1 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=0.1116p ps=0.98u w=0.36u l=0.5u
X2411 a_8064_5176 a_7652_4855 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2412 a_12068_5644 a_10900_6040 a_11864_5644 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2413 vccd1 a_6558_7080 a_6426_7124 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2414 a_33440_6428 a_22560_4292 vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=0.2016p ps=1.48u w=0.36u l=0.6u
X2415 a_8277_6916 a_8157_6296 a_7533_6296 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2416 SDAC[7] a_32236_3160 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2417 a_16271_5557 a_6252_7864 vccd1 vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.3718p ps=2.57u w=0.845u l=0.5u
X2418 vssd1 a_24675_4728 a_23320_6574 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2419 vssd1 a_5129_4336 a_5024_4476 vssd1 nfet_06v0 ad=0.1224p pd=1.04u as=94.5f ps=0.885u w=0.36u l=0.6u
X2420 SC a_35708_9001 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2421 a_15324_6608 a_21392_8392 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2422 vccd1 a_35916_7168 a_35812_7212 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2423 a_31100_9831 a_30792_9880 vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X2424 a_23052_7564 a_24435_7098 a_25367_7608 vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2425 vccd1 a_3932_9783 a_3844_9880 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2426 a_5948_11784 a_5860_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2427 vssd1 a_28757_3989 a_29044_12359 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2428 a_13656_7212 a_13104_7195 a_13452_7212 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2429 a_25718_12404 a_25242_11828 vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2430 a_31561_4336 a_22560_4292 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
D121 a_2468_3254 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2431 vssd1 a_9408_3608 SDAC[0] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2432 a_23616_4476 a_21092_4472 a_23304_4476 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2433 a_11508_8780 a_10340_9176 a_11304_8780 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2434 vccd1 a_24872_6428 a_25289_6384 vccd1 pfet_06v0 ad=0.44p pd=2.88u as=0.26p ps=1.52u w=1u l=0.5u
X2435 a_7486_7124 a_7050_7124 a_7254_7124 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2436 SDAC[4] a_21504_3608 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2437 a_30613_8462 a_30493_7864 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X2438 a_30613_5326 a_30493_4728 vccd1 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.379p ps=2.37u w=0.36u l=0.5u
X2439 vssd1 a_22560_4292 a_28336_6044 vssd1 nfet_06v0 ad=0.2016p pd=1.48u as=43.199997f ps=0.6u w=0.36u l=0.6u
D122 a_1908_4118 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2440 vssd1 a_26902_12404 a_27378_12403 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X2441 vccd1 a_22364_4032 a_22260_4076 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2442 a_23599_5996 a_23721_4336 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2443 a_19797_9477 a_18793_9520 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2444 a_18244_7124 a_17640_7564 vccd1 vccd1 pfet_06v0 ad=0.1456p pd=1.08u as=0.4005p ps=2.12u w=0.56u l=0.5u
X2445 vccd1 a_28540_9500 a_26456_8736 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2446 a_24360_9152 a_19524_11448 vssd1 vssd1 nfet_06v0 ad=0.1584p pd=1.6u as=0.153p ps=1.195u w=0.36u l=0.6u
X2447 vccd1 a_3564_7864 a_1772_7864 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2448 vccd1 a_20495_6296 a_21871_5250 vccd1 pfet_06v0 ad=0.2197p pd=1.365u as=0.2197p ps=1.365u w=0.845u l=0.5u
X2449 vssd1 a_15324_6608 a_13496_6366 vssd1 nfet_06v0 ad=0.1053p pd=0.925u as=0.1782p ps=1.69u w=0.405u l=0.6u
X2450 vccd1 a_24976_3608 SDAC[5] vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2451 a_19297_6341 a_15483_8723 vssd1 vssd1 nfet_06v0 ad=0.1304p pd=1.135u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2452 a_6558_7080 a_5689_5904 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2453 a_20060_11784 a_19972_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2454 vssd1 a_19052_8648 a_18760_8692 vssd1 nfet_06v0 ad=0.218p pd=1.52u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2455 a_8820_5176 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
X2456 vssd1 a_15568_5176 SDAC[2] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2457 vssd1 a_35737_5996 a_35668_6044 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=62.1f ps=0.705u w=0.36u l=0.6u
X2458 a_11660_5644 a_11560_5600 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X2459 a_27216_9180 a_27068_8736 a_27048_9180 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=43.199997f ps=0.6u w=0.36u l=0.6u
X2460 a_29128_6044 a_27328_5627 a_28188_5600 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2461 a_9868_6744 a_9768_6574 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2462 a_37500_4728 a_37108_11089 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4015p ps=1.92u w=1.22u l=0.5u
X2463 a_4488_7612 a_2276_7608 a_3548_7168 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X2464 vssd1 a_6440_9152 a_3564_7864 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X2465 vccd1 a_35708_9001 SC vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2466 a_23599_5996 a_23721_4336 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2467 vssd1 a_12556_4773 a_12468_4817 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2468 a_22660_5176 a_22932_4728 a_22848_5176 vccd1 pfet_06v0 ad=0.44955p pd=1.955u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2469 a_14280_9152 a_14540_8648 vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X2470 a_22748_10216 a_22660_10260 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2471 vccd1 a_21180_4416 a_25124_4472 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2472 a_33094_5892 a_31465_5512 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.4941p ps=2.03u w=1.22u l=0.5u
X2473 a_6558_7080 a_5689_5904 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2474 a_16257_4476 a_1908_4118 vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X2475 a_37396_5176 a_36972_7864 a_37152_5194 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4248p ps=1.94u w=1.22u l=0.5u
X2476 a_25312_5556 a_5972_3608 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2477 a_6133_8693 a_5129_9040 vccd1 vccd1 pfet_06v0 ad=0.5346p pd=3.31u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2478 vccd1 a_21392_8392 a_15324_6608 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2479 SDAC[1] a_13216_3608 vssd1 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2480 a_31117_7864 a_31509_7864 vssd1 vssd1 nfet_06v0 ad=0.333p pd=2.57u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2481 a_11100_8780 a_11000_8736 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X2482 a_5024_4476 a_2500_4472 a_4712_4476 vssd1 nfet_06v0 ad=94.5f pd=0.885u as=0.2007p ps=1.475u w=0.36u l=0.6u
X2483 a_21628_11784 a_21540_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2484 vccd1 a_21180_4416 a_22660_6423 vccd1 pfet_06v0 ad=0.2249p pd=1.385u as=0.3806p ps=2.61u w=0.865u l=0.5u
X2485 a_11737_6384 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.26p pd=1.52u as=0.29465p ps=1.74u w=1u l=0.5u
X2486 vccd1 a_10035_7080 a_9903_7124 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2487 SDAC[6] a_28428_3160 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
D123 vssd1 a_1908_4118 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2488 a_21356_8736 a_21048_8780 vssd1 vssd1 nfet_06v0 ad=0.2007p pd=1.475u as=0.2016p ps=1.48u w=0.36u l=0.6u
X2489 a_34832_5627 a_34420_6040 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2490 vssd1 a_30499_10653 a_28540_9500 vssd1 nfet_06v0 ad=0.282625p pd=1.87u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2491 SDAC[7] a_32236_3160 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.5368p ps=3.32u w=1.22u l=0.5u
X2492 vccd1 a_22560_4292 a_34364_5176 vccd1 pfet_06v0 ad=0.45p pd=2.02u as=0.3432p ps=2.44u w=0.78u l=0.5u
X2493 a_26734_12404 a_26070_11828 vssd1 vssd1 nfet_06v0 ad=43.199997f pd=0.6u as=93.59999f ps=0.88u w=0.36u l=0.6u
X2494 vssd1 a_18236_7864 a_18172_7908 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.1312p ps=1.14u w=0.82u l=0.6u
X2495 vccd1 a_31453_10792 a_31573_10260 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2496 a_25374_11784 a_37513_5984 vssd1 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.3586p ps=2.51u w=0.815u l=0.6u
X2497 a_14616_9477 a_14876_9477 vccd1 vccd1 pfet_06v0 ad=0.462p pd=2.98u as=0.4015p ps=1.92u w=1.05u l=0.5u
X2498 a_25884_4076 a_25784_4032 vssd1 vssd1 nfet_06v0 ad=93.59999f pd=0.88u as=0.1584p ps=1.6u w=0.36u l=0.6u
X2499 a_4145_3608 a_2468_3254 vccd1 vccd1 pfet_06v0 ad=0.2938p pd=1.65u as=0.4972p ps=3.14u w=1.13u l=0.5u
D124 a_2468_4822 vccd1 diode_pd2nw_06v0 pj=1.86u area=0.2052p
X2500 a_4800_7612 a_2688_7195 a_4488_7612 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X2501 vccd1 a_2588_9783 a_2500_9880 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2502 a_21504_4059 a_21092_4472 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2503 SDAC[2] a_15568_5176 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2504 a_18376_9564 a_16164_9559 a_17436_9831 vccd1 pfet_06v0 ad=0.25375p pd=1.51u as=0.2424p ps=1.465u w=0.505u l=0.5u
X2505 vccd1 a_6496_3988 a_1908_4118 vccd1 pfet_06v0 ad=0.3172p pd=1.74u as=0.4392p ps=1.94u w=1.22u l=0.5u
X2506 vccd1 a_2588_6647 a_2500_6744 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2507 a_6508_11351 a_6420_11448 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2508 a_35812_7212 a_1908_4118 vccd1 vccd1 pfet_06v0 ad=0.3432p pd=2.44u as=0.45p ps=2.02u w=0.78u l=0.5u
D125 vssd1 a_2916_4822 diode_nd2ps_06v0 pj=1.86u area=0.2052p
X2509 a_27028_6340 a_23756_7080 a_27236_6340 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2510 a_34144_9238 a_34292_8648 a_34144_8693 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.44955p ps=1.955u w=1.215u l=0.5u
X2511 SDAC[5] a_24976_3608 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2512 vssd1 a_24976_3608 SDAC[5] vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2513 a_9892_6040 a_2468_4822 a_7416_8142 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2514 a_3472_5627 a_3060_6040 vssd1 vssd1 nfet_06v0 ad=0.1782p pd=1.69u as=0.1053p ps=0.925u w=0.405u l=0.6u
X2515 a_8086_7700 a_7254_7124 a_7938_7124 vccd1 pfet_06v0 ad=0.3852p pd=2.86u as=61.199993f ps=0.7u w=0.36u l=0.5u
X2516 a_30700_11784 a_30612_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2517 a_27609_11448 a_26879_11044 vccd1 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
X2518 a_31100_9831 a_30792_9880 vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X2519 a_15324_6608 a_21392_8392 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X2520 a_3464_4076 a_2912_4059 a_3260_4076 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2521 vssd1 a_23599_5996 a_23535_6040 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2522 vssd1 a_25248_9120 a_24876_3160 vssd1 nfet_06v0 ad=0.2344p pd=1.56u as=0.3608p ps=2.52u w=0.82u l=0.6u
X2523 a_34441_11828 a_33711_11850 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.282625p ps=1.87u w=0.82u l=0.6u
X2524 vssd1 a_11279_7864 a_11215_7909 vssd1 nfet_06v0 ad=0.3586p pd=2.51u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2525 a_17418_6916 a_17318_6562 a_16694_6296 vccd1 pfet_06v0 ad=61.199993f pd=0.7u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2526 vccd1 a_26163_11000 a_26031_11044 vccd1 pfet_06v0 ad=0.1116p pd=0.98u as=0.3852p ps=2.86u w=0.36u l=0.5u
X2527 a_12860_7909 a_16271_5557 a_16833_7909 vssd1 nfet_06v0 ad=0.2119p pd=1.335u as=0.1304p ps=1.135u w=0.815u l=0.6u
X2528 COMP_CLK a_33916_11000 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2529 vssd1 a_35708_11000 a_33916_11000 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2530 a_37168_10748 a_35056_10331 a_36856_10748 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X2531 a_28428_3160 a_30220_3160 vccd1 vccd1 pfet_06v0 ad=0.3782p pd=1.84u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2532 a_35232_4860 a_33511_5187 a_34104_5118 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2533 a_31844_6040 a_2468_4822 a_31509_7864 vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2534 a_28801_9180 a_1908_4118 vssd1 vssd1 nfet_06v0 ad=0.134p pd=1.1u as=0.1224p ps=1.04u w=0.36u l=0.6u
X2535 vccd1 a_30924_11351 a_30836_11448 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.5368p ps=3.32u w=1.22u l=1u
X2536 vssd1 a_34441_11828 a_36268_12281 vssd1 nfet_06v0 ad=0.2244p pd=1.9u as=0.2569p ps=1.56u w=0.51u l=0.6u
X2537 a_36833_6044 a_22560_4292 vccd1 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.3432p ps=2.44u w=0.78u l=0.5u
X2538 a_34000_6428 a_32279_6755 a_32872_6686 vccd1 pfet_06v0 ad=0.2028p pd=1.3u as=0.2028p ps=1.3u w=0.78u l=0.5u
X2539 vssd1 a_9408_3608 SDAC[0] vssd1 nfet_06v0 ad=0.2132p pd=1.34u as=0.2132p ps=1.34u w=0.82u l=0.6u
X2540 a_8636_11784 a_8548_11828 vssd1 vssd1 nfet_06v0 ad=0.3608p pd=2.52u as=0.3608p ps=2.52u w=0.82u l=1u
X2541 vccd1 a_24115_5557 a_26804_7953 vccd1 pfet_06v0 ad=0.4015p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X2542 a_18688_9564 a_16576_9880 a_18376_9564 vccd1 pfet_06v0 ad=0.1313p pd=1.025u as=0.25375p ps=1.51u w=0.505u l=0.5u
X2543 a_8028_8263 a_7720_8312 vccd1 vccd1 pfet_06v0 ad=0.2424p pd=1.465u as=0.2222p ps=1.89u w=0.505u l=0.5u
X2544 vccd1 a_35708_11000 a_33916_11000 vccd1 pfet_06v0 ad=0.5368p pd=3.32u as=0.3782p ps=1.84u w=1.22u l=0.5u
X2545 vssd1 a_37912_11045 a_35708_11000 vssd1 nfet_06v0 ad=0.153p pd=1.195u as=0.2178p ps=1.87u w=0.495u l=0.6u
X2546 vccd1 a_2916_4822 a_7799_5557 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.3159p ps=1.735u w=1.215u l=0.5u
X2547 a_23107_5557 a_20028_7080 a_22919_5557 vccd1 pfet_06v0 ad=0.3159p pd=1.735u as=0.5346p ps=3.31u w=1.215u l=0.5u
X2548 a_21891_4772 a_6252_7864 vssd1 vssd1 nfet_06v0 ad=0.1517p pd=1.19u as=0.3608p ps=2.52u w=0.82u l=0.6u
.ends

