* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt TOP top_c5 top_c3 top_c2 top_c4 top_c0 top_c1 top_c_dummy common_bottom
X0 top_c5.t0 common_bottom.t39 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X1 top_c3.t0 common_bottom.t55 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X2 top_c5.t1 common_bottom.t38 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X3 top_c3.t1 common_bottom.t3 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X4 top_c4.t0 common_bottom.t44 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X5 top_c5.t2 common_bottom.t37 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X6 top_c5.t3 common_bottom.t36 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X7 top_c5.t4 common_bottom.t35 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X8 top_c5.t5 common_bottom.t34 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X9 top_c0.t0 common_bottom.t57 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X10 top_c5.t6 common_bottom.t33 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X11 top_c3.t2 common_bottom.t7 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X12 top_c5.t7 common_bottom.t32 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X13 top_c3.t3 common_bottom.t54 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X14 top_c5.t8 common_bottom.t31 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X15 top_c5.t9 common_bottom.t30 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X16 top_c2.t0 common_bottom.t49 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X17 top_c5.t10 common_bottom.t29 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X18 top_c4.t1 common_bottom.t2 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X19 top_c3.t4 common_bottom.t62 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X20 top_c4.t2 common_bottom.t60 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X21 top_c5.t11 common_bottom.t28 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X22 top_c5.t12 common_bottom.t27 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X23 top_c5.t13 common_bottom.t26 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X24 top_c4.t3 common_bottom.t47 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X25 top_c4.t4 common_bottom.t6 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X26 top_c4.t5 common_bottom.t41 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X27 top_c5.t14 common_bottom.t25 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X28 top_c5.t15 common_bottom.t24 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X29 top_c4.t6 common_bottom.t43 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X30 top_c4.t7 common_bottom.t1 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X31 top_c5.t16 common_bottom.t23 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X32 top_c5.t17 common_bottom.t22 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X33 top_c5.t18 common_bottom.t21 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X34 top_c4.t8 common_bottom.t46 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X35 top_c2.t1 common_bottom.t63 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X36 top_c4.t9 common_bottom.t5 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X37 top_c5.t19 common_bottom.t20 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X38 top_c_dummy.t0 common_bottom.t58 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X39 top_c5.t20 common_bottom.t19 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X40 top_c2.t2 common_bottom.t52 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X41 top_c5.t21 common_bottom.t18 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X42 top_c0.t1 common_bottom.t59 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X43 top_c5.t22 common_bottom.t17 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X44 top_c4.t10 common_bottom.t40 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X45 top_c5.t23 common_bottom.t16 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X46 top_c1.t0 common_bottom.t4 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X47 top_c5.t24 common_bottom.t15 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X48 top_c4.t11 common_bottom.t42 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X49 top_c4.t12 common_bottom.t0 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X50 top_c5.t25 common_bottom.t14 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X51 top_c3.t5 common_bottom.t56 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X52 top_c4.t13 common_bottom.t50 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X53 top_c4.t14 common_bottom.t48 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X54 top_c5.t26 common_bottom.t13 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X55 top_c5.t27 common_bottom.t12 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X56 top_c3.t6 common_bottom.t61 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X57 top_c4.t15 common_bottom.t51 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X58 top_c5.t28 common_bottom.t11 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X59 top_c5.t29 common_bottom.t10 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X60 top_c5.t30 common_bottom.t9 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X61 top_c3.t7 common_bottom.t53 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X62 top_c2.t3 common_bottom.t45 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
X63 top_c5.t31 common_bottom.t8 cap_mim_2f0_m4m5_noshield c_width=7u c_length=7u
R0 top_c5.n59 top_c5.n58 47.7486
R1 top_c5.n26 top_c5.n9 10.9483
R2 top_c5.n58 top_c5.n47 6.64428
R3 top_c5.n47 top_c5.n46 5.79894
R4 top_c5.n58 top_c5.n57 4.31368
R5 top_c5.n47 top_c5.n29 4.28582
R6 top_c5.n27 top_c5.n1 4.28582
R7 top_c5.n28 top_c5.n0 4.28582
R8 top_c5.n26 top_c5.n25 4.27886
R9 top_c5.n28 top_c5.n27 3.26928
R10 top_c5.n27 top_c5.n26 3.26768
R11 top_c5.n59 top_c5.n28 2.51351
R12 top_c5.n51 top_c5.n49 0.988357
R13 top_c5.n49 top_c5.n48 0.988357
R14 top_c5.n36 top_c5.n35 0.988357
R15 top_c5.n38 top_c5.n35 0.988357
R16 top_c5.n41 top_c5.n34 0.988357
R17 top_c5.n12 top_c5.n11 0.988357
R18 top_c5.n14 top_c5.n11 0.988357
R19 top_c5.n17 top_c5.n10 0.988357
R20 top_c5.n19 top_c5.n10 0.988357
R21 top_c5.n24 top_c5.n23 0.988357
R22 top_c5.n3 top_c5.n2 0.988357
R23 top_c5.n5 top_c5.n3 0.988357
R24 top_c5.n43 top_c5.n34 0.988261
R25 top_c5.n33 top_c5.n32 0.987576
R26 top_c5.n44 top_c5.n33 0.960525
R27 top_c5.n56 top_c5.n48 0.9605
R28 top_c5.n54 top_c5.n51 0.9605
R29 top_c5.n30 top_c5.n29 0.9605
R30 top_c5.n1 top_c5.n0 0.9605
R31 top_c5.n23 top_c5.n21 0.9605
R32 top_c5.n6 top_c5.n5 0.9605
R33 top_c5.n8 top_c5.n2 0.9605
R34 top_c5.n25 top_c5.n1 0.9575
R35 top_c5.n36 top_c5.t2 0.60448
R36 top_c5.n12 top_c5.t5 0.60448
R37 top_c5.n6 top_c5.t18 0.60448
R38 top_c5.n46 top_c5.n45 0.59544
R39 top_c5.n52 top_c5.t25 0.586765
R40 top_c5.n40 top_c5.n39 0.5405
R41 top_c5.n16 top_c5.n15 0.5405
R42 top_c5.n53 top_c5.n52 0.526689
R43 top_c5.n54 top_c5.n53 0.512643
R44 top_c5.n41 top_c5.n40 0.512643
R45 top_c5.n17 top_c5.n16 0.512643
R46 top_c5.n57 top_c5.n56 0.512643
R47 top_c5.n39 top_c5.n38 0.512643
R48 top_c5.n15 top_c5.n14 0.512643
R49 top_c5.n9 top_c5.n8 0.512643
R50 top_c5 top_c5.n59 0.494375
R51 top_c5.n44 top_c5.n43 0.484786
R52 top_c5.n21 top_c5.n19 0.484786
R53 top_c5.n46 top_c5.n30 0.322414
R54 top_c5.n52 top_c5.t10 0.106765
R55 top_c5.n53 top_c5.t23 0.0923367
R56 top_c5.n49 top_c5.t11 0.0923367
R57 top_c5.n50 top_c5.t26 0.0923367
R58 top_c5.n55 top_c5.t12 0.0923367
R59 top_c5.n57 top_c5.t29 0.0923367
R60 top_c5.n35 top_c5.t8 0.0923367
R61 top_c5.n37 top_c5.t24 0.0923367
R62 top_c5.n39 top_c5.t13 0.0923367
R63 top_c5.n40 top_c5.t27 0.0923367
R64 top_c5.n34 top_c5.t28 0.0923367
R65 top_c5.n42 top_c5.t14 0.0923367
R66 top_c5.n32 top_c5.t30 0.0923367
R67 top_c5.n31 top_c5.t16 0.0923367
R68 top_c5.n45 top_c5.t0 0.0923367
R69 top_c5.n11 top_c5.t7 0.0923367
R70 top_c5.n13 top_c5.t22 0.0923367
R71 top_c5.n15 top_c5.t1 0.0923367
R72 top_c5.n16 top_c5.t15 0.0923367
R73 top_c5.n10 top_c5.t31 0.0923367
R74 top_c5.n18 top_c5.t17 0.0923367
R75 top_c5.n20 top_c5.t4 0.0923367
R76 top_c5.n22 top_c5.t20 0.0923367
R77 top_c5.n24 top_c5.t6 0.0923367
R78 top_c5.n3 top_c5.t21 0.0923367
R79 top_c5.n4 top_c5.t3 0.0923367
R80 top_c5.n7 top_c5.t19 0.0923367
R81 top_c5.n9 top_c5.t9 0.0923367
R82 top_c5.n25 top_c5.n24 0.0293187
R83 top_c5.n33 top_c5.n31 0.029221
R84 top_c5.n50 top_c5.n48 0.0283571
R85 top_c5.n51 top_c5.n50 0.0283571
R86 top_c5.n56 top_c5.n55 0.0283571
R87 top_c5.n55 top_c5.n54 0.0283571
R88 top_c5.n38 top_c5.n37 0.0283571
R89 top_c5.n37 top_c5.n36 0.0283571
R90 top_c5.n43 top_c5.n42 0.0283571
R91 top_c5.n42 top_c5.n41 0.0283571
R92 top_c5.n32 top_c5.n29 0.0283571
R93 top_c5.n31 top_c5.n30 0.0283571
R94 top_c5.n45 top_c5.n44 0.0283571
R95 top_c5.n13 top_c5.n12 0.0283571
R96 top_c5.n14 top_c5.n13 0.0283571
R97 top_c5.n18 top_c5.n17 0.0283571
R98 top_c5.n19 top_c5.n18 0.0283571
R99 top_c5.n21 top_c5.n20 0.0283571
R100 top_c5.n20 top_c5.n0 0.0283571
R101 top_c5.n23 top_c5.n22 0.0283571
R102 top_c5.n22 top_c5.n1 0.0283571
R103 top_c5.n5 top_c5.n4 0.0283571
R104 top_c5.n4 top_c5.n2 0.0283571
R105 top_c5.n7 top_c5.n6 0.0283571
R106 top_c5.n8 top_c5.n7 0.0283571
R107 common_bottom common_bottom.t6 6.59189
R108 common_bottom.t50 common_bottom.t54 1.23983
R109 common_bottom.t54 common_bottom.t37 1.23983
R110 common_bottom.t37 common_bottom.t15 1.23983
R111 common_bottom.t15 common_bottom.t26 1.23983
R112 common_bottom.t12 common_bottom.t26 1.23983
R113 common_bottom.t25 common_bottom.t12 1.23983
R114 common_bottom.t56 common_bottom.t34 1.23216
R115 common_bottom.t52 common_bottom.t28 1.23216
R116 common_bottom.t13 common_bottom.t7 1.23216
R117 common_bottom.t27 common_bottom.t16 1.23216
R118 common_bottom.t61 common_bottom.t49 1.23216
R119 common_bottom.t47 common_bottom.t0 1.23216
R120 common_bottom.t62 common_bottom.t11 1.23216
R121 common_bottom.t34 common_bottom.t17 1.23216
R122 common_bottom.t17 common_bottom.t38 1.23216
R123 common_bottom.t32 common_bottom.t5 1.23216
R124 common_bottom.t4 common_bottom.t44 1.23216
R125 common_bottom.t29 common_bottom.t58 1.23216
R126 common_bottom.t14 common_bottom.t57 1.23216
R127 common_bottom.t48 common_bottom.t31 1.23216
R128 common_bottom.t31 common_bottom.t63 1.23216
R129 common_bottom.t24 common_bottom.t22 1.23216
R130 common_bottom.t22 common_bottom.t35 1.23216
R131 common_bottom.t19 common_bottom.t8 1.23216
R132 common_bottom.t33 common_bottom.t46 1.23216
R133 common_bottom.t40 common_bottom.t3 1.23216
R134 common_bottom.t30 common_bottom.t20 1.23216
R135 common_bottom.t42 common_bottom.t36 1.23216
R136 common_bottom.t2 common_bottom.t18 1.23216
R137 common_bottom.t39 common_bottom.t25 1.23216
R138 common_bottom.t56 common_bottom.t28 1.2245
R139 common_bottom.t13 common_bottom.t28 1.2245
R140 common_bottom.t13 common_bottom.t27 1.2245
R141 common_bottom.t27 common_bottom.t61 1.2245
R142 common_bottom.t61 common_bottom.t47 1.2245
R143 common_bottom.t11 common_bottom.t47 1.2245
R144 common_bottom.t11 common_bottom.t25 1.2245
R145 common_bottom.t5 common_bottom.t38 1.2245
R146 common_bottom.t44 common_bottom.t5 1.2245
R147 common_bottom.t58 common_bottom.t44 1.2245
R148 common_bottom.t57 common_bottom.t58 1.2245
R149 common_bottom.t59 common_bottom.t57 1.2245
R150 common_bottom.t62 common_bottom.t12 1.2245
R151 common_bottom.t62 common_bottom.t0 1.2245
R152 common_bottom.t0 common_bottom.t49 1.2245
R153 common_bottom.t49 common_bottom.t16 1.2245
R154 common_bottom.t16 common_bottom.t7 1.2245
R155 common_bottom.t7 common_bottom.t52 1.2245
R156 common_bottom.t34 common_bottom.t52 1.2245
R157 common_bottom.t17 common_bottom.t32 1.2245
R158 common_bottom.t32 common_bottom.t52 1.2245
R159 common_bottom.t32 common_bottom.t4 1.2245
R160 common_bottom.t4 common_bottom.t7 1.2245
R161 common_bottom.t4 common_bottom.t29 1.2245
R162 common_bottom.t29 common_bottom.t16 1.2245
R163 common_bottom.t29 common_bottom.t14 1.2245
R164 common_bottom.t14 common_bottom.t49 1.2245
R165 common_bottom.t60 common_bottom.t59 1.2245
R166 common_bottom.t14 common_bottom.t60 1.2245
R167 common_bottom.t60 common_bottom.t0 1.2245
R168 common_bottom.t48 common_bottom.t26 1.2245
R169 common_bottom.t60 common_bottom.t48 1.2245
R170 common_bottom.t48 common_bottom.t62 1.2245
R171 common_bottom.t31 common_bottom.t15 1.2245
R172 common_bottom.t31 common_bottom.t59 1.2245
R173 common_bottom.t63 common_bottom.t37 1.2245
R174 common_bottom.t63 common_bottom.t55 1.2245
R175 common_bottom.t55 common_bottom.t59 1.2245
R176 common_bottom.t55 common_bottom.t21 1.2245
R177 common_bottom.t21 common_bottom.t57 1.2245
R178 common_bottom.t21 common_bottom.t45 1.2245
R179 common_bottom.t45 common_bottom.t3 1.2245
R180 common_bottom.t45 common_bottom.t58 1.2245
R181 common_bottom.t45 common_bottom.t1 1.2245
R182 common_bottom.t1 common_bottom.t44 1.2245
R183 common_bottom.t1 common_bottom.t53 1.2245
R184 common_bottom.t53 common_bottom.t5 1.2245
R185 common_bottom.t53 common_bottom.t24 1.2245
R186 common_bottom.t24 common_bottom.t38 1.2245
R187 common_bottom.t35 common_bottom.t19 1.2245
R188 common_bottom.t22 common_bottom.t8 1.2245
R189 common_bottom.t53 common_bottom.t8 1.2245
R190 common_bottom.t46 common_bottom.t3 1.2245
R191 common_bottom.t8 common_bottom.t46 1.2245
R192 common_bottom.t1 common_bottom.t46 1.2245
R193 common_bottom.t19 common_bottom.t33 1.2245
R194 common_bottom.t33 common_bottom.t40 1.2245
R195 common_bottom.t30 common_bottom.t42 1.2245
R196 common_bottom.t40 common_bottom.t30 1.2245
R197 common_bottom.t3 common_bottom.t20 1.2245
R198 common_bottom.t21 common_bottom.t20 1.2245
R199 common_bottom.t20 common_bottom.t36 1.2245
R200 common_bottom.t55 common_bottom.t36 1.2245
R201 common_bottom.t54 common_bottom.t18 1.2245
R202 common_bottom.t36 common_bottom.t18 1.2245
R203 common_bottom.t63 common_bottom.t18 1.2245
R204 common_bottom.t42 common_bottom.t2 1.2245
R205 common_bottom.t2 common_bottom.t50 1.2245
R206 common_bottom.t23 common_bottom.t39 1.2245
R207 common_bottom.t11 common_bottom.t23 1.2245
R208 common_bottom.t23 common_bottom.t9 1.2245
R209 common_bottom.t9 common_bottom.t47 1.2245
R210 common_bottom.t9 common_bottom.t43 1.2245
R211 common_bottom.t43 common_bottom.t61 1.2245
R212 common_bottom.t43 common_bottom.t10 1.2245
R213 common_bottom.t10 common_bottom.t27 1.2245
R214 common_bottom.t10 common_bottom.t41 1.2245
R215 common_bottom.t41 common_bottom.t13 1.2245
R216 common_bottom.t41 common_bottom.t51 1.2245
R217 common_bottom.t28 common_bottom.t51 1.2245
R218 common_bottom.t6 common_bottom.t51 1.2245
R219 common_bottom.t6 common_bottom.t56 1.2245
R220 top_c3.n6 top_c3.n5 24.4226
R221 top_c3.n3 top_c3.t4 11.0947
R222 top_c3.n0 top_c3.t3 11.0893
R223 top_c3.n1 top_c3.n0 6.64802
R224 top_c3.n2 top_c3.n1 6.64673
R225 top_c3.n4 top_c3.n3 6.64471
R226 top_c3.n5 top_c3.n4 6.64471
R227 top_c3.n6 top_c3.n2 5.28193
R228 top_c3.n0 top_c3.t0 4.60328
R229 top_c3.n2 top_c3.t7 4.6016
R230 top_c3.n3 top_c3.t6 4.59742
R231 top_c3.n5 top_c3.t5 4.59742
R232 top_c3.n4 top_c3.t2 4.45045
R233 top_c3.n1 top_c3.t1 4.44401
R234 top_c3 top_c3.n6 1.0805
R235 top_c4.n28 top_c4.n27 31.4494
R236 top_c4.n21 top_c4.n20 9.65716
R237 top_c4.n22 top_c4.n15 9.6293
R238 top_c4.n23 top_c4.n14 9.6293
R239 top_c4.n26 top_c4.n25 9.6293
R240 top_c4.n7 top_c4.n6 9.36076
R241 top_c4.n4 top_c4.n1 9.3329
R242 top_c4.n5 top_c4.n0 9.3329
R243 top_c4.n28 top_c4.n12 8.94299
R244 top_c4.n19 top_c4.n18 7.62953
R245 top_c4.n20 top_c4.n19 5.96827
R246 top_c4.n8 top_c4.n7 5.96198
R247 top_c4.n2 top_c4.n1 5.32736
R248 top_c4.n19 top_c4.t6 4.58128
R249 top_c4.n12 top_c4.n11 4.50243
R250 top_c4.n27 top_c4.n13 4.49219
R251 top_c4.n8 top_c4.t10 4.43431
R252 top_c4.n12 top_c4.n8 3.27471
R253 top_c4.n27 top_c4.n26 2.59314
R254 top_c4.n15 top_c4.n14 1.913
R255 top_c4.n1 top_c4.n0 1.913
R256 top_c4.n20 top_c4.n15 1.463
R257 top_c4.n26 top_c4.n14 1.463
R258 top_c4.n7 top_c4.n0 1.463
R259 top_c4 top_c4.n28 0.8105
R260 top_c4.n16 top_c4.t14 0.586765
R261 top_c4.n9 top_c4.t9 0.586765
R262 top_c4.n18 top_c4.n17 0.5405
R263 top_c4.n11 top_c4.n10 0.5405
R264 top_c4.n17 top_c4.n16 0.526689
R265 top_c4.n10 top_c4.n9 0.526689
R266 top_c4.n23 top_c4.n22 0.484786
R267 top_c4.n5 top_c4.n4 0.484786
R268 top_c4.n25 top_c4.n13 0.482942
R269 top_c4.n2 top_c4.t13 0.307092
R270 top_c4.n3 top_c4.n2 0.297766
R271 top_c4.n13 top_c4.t4 0.113497
R272 top_c4.n16 top_c4.t2 0.106765
R273 top_c4.n9 top_c4.t0 0.106765
R274 top_c4.n24 top_c4.t15 0.0923367
R275 top_c4.n21 top_c4.t5 0.0923367
R276 top_c4.n17 top_c4.t12 0.0923367
R277 top_c4.n18 top_c4.t3 0.0923367
R278 top_c4.n10 top_c4.t7 0.0923367
R279 top_c4.n11 top_c4.t8 0.0923367
R280 top_c4.n6 top_c4.t11 0.0923367
R281 top_c4.n3 top_c4.t1 0.0923367
R282 top_c4.n24 top_c4.n23 0.0283571
R283 top_c4.n25 top_c4.n24 0.0283571
R284 top_c4.n22 top_c4.n21 0.0283571
R285 top_c4.n6 top_c4.n5 0.0283571
R286 top_c4.n4 top_c4.n3 0.0283571
R287 top_c0 top_c0.n0 16.4389
R288 top_c0.n0 top_c0.t1 7.71362
R289 top_c0.n0 top_c0.t0 4.44401
R290 top_c2.n2 top_c2.n1 21.2892
R291 top_c2.n1 top_c2.t0 14.4679
R292 top_c2.n0 top_c2.t1 14.4636
R293 top_c2.n2 top_c2.n0 11.7153
R294 top_c2.n1 top_c2.t2 4.45022
R295 top_c2.n0 top_c2.t3 4.44401
R296 top_c2 top_c2.n2 1.37413
R297 top_c_dummy top_c_dummy.t0 17.5392
R298 top_c1 top_c1.t0 14.1391
C0 top_c3 top_c_dummy 0.084329f
C1 top_c3 top_c2 2.97689f
C2 top_c0 top_c1 3.2923f
C3 top_c4 m3_13080_37400 0.177159f
C4 top_c_dummy top_c5 0.619868f
C5 top_c4 m3_9610_37600 0.290507f
C6 top_c1 top_c4 0.448342f
C7 top_c2 top_c5 2.21258f
C8 common_bottom m3_n1905_37400 0.979483f
C9 top_c0 top_c_dummy 0.554286f
C10 top_c1 m3_9610_37600 0.135476f
C11 top_c0 top_c2 0.090243f
C12 m3_1090_37400 top_c2 0.27095f
C13 top_c4 top_c_dummy 0.491368f
C14 common_bottom top_c3 10.3733f
C15 top_c3 m3_n1905_37400 0.245343f
C16 top_c4 top_c2 0.740292f
C17 top_c2 m3_13080_37400 0.029917f
C18 common_bottom top_c5 32.068798f
C19 top_c5 m3_n1905_37400 0.720308f
C20 top_c1 top_c_dummy 0.013558f
C21 top_c2 m3_9610_37600 3.18752f
C22 common_bottom m3_16090_37400 0.97451f
C23 top_c1 top_c2 0.077876f
C24 top_c3 top_c5 2.96266f
C25 common_bottom top_c0 3.10669f
C26 common_bottom m3_1090_37400 0.975713f
C27 top_c3 m3_16090_37400 0.018825f
C28 common_bottom top_c4 17.471699f
C29 top_c4 m3_n1905_37400 3.33663f
C30 top_c2 top_c_dummy 3.46169f
C31 top_c0 top_c3 0.200626f
C32 m3_16090_37400 top_c5 0.592178f
C33 common_bottom m3_13080_37400 1.11323f
C34 top_c3 m3_1090_37400 3.38043f
C35 common_bottom m3_9610_37600 0.974327f
C36 top_c3 top_c4 4.93972f
C37 common_bottom top_c1 2.03298f
C38 top_c0 top_c5 0.88364f
C39 m3_1090_37400 top_c5 0.434547f
C40 top_c3 m3_13080_37400 3.57081f
C41 top_c4 top_c5 8.98776f
C42 top_c3 m3_9610_37600 0.026795f
C43 top_c1 top_c3 0.200621f
C44 top_c4 m3_16090_37400 3.74506f
C45 common_bottom top_c_dummy 2.01547f
C46 top_c5 m3_13080_37400 0.805341f
C47 common_bottom top_c2 6.66733f
C48 m3_9610_37600 top_c5 0.683089f
C49 top_c0 top_c4 0.448241f
C50 top_c1 top_c5 1.04224f
C51 top_c4 m3_1090_37400 0.152828f
C52 common_bottom VSUBS 81.92847f
C53 top_c1 VSUBS 7.456892f
C54 top_c0 VSUBS 9.766644f
C55 top_c_dummy VSUBS 8.100149f
C56 top_c2 VSUBS 19.239426f
C57 top_c3 VSUBS 28.22961f
C58 top_c4 VSUBS 44.97781f
C59 top_c5 VSUBS 85.22208f
C60 m3_16090_37400 VSUBS 4.75247f $ **FLOATING
C61 m3_13080_37400 VSUBS 4.85576f $ **FLOATING
C62 m3_9610_37600 VSUBS 4.70657f $ **FLOATING
C63 m3_1090_37400 VSUBS 4.78423f $ **FLOATING
C64 m3_n1905_37400 VSUBS 4.76133f $ **FLOATING
C65 top_c1.t0 VSUBS 5.10351f
C66 top_c_dummy.t0 VSUBS 4.65036f
C67 top_c2.t1 VSUBS 4.29711f
C68 top_c2.t3 VSUBS 3.78188f
C69 top_c2.n0 VSUBS 1.10189f
C70 top_c2.t0 VSUBS 3.68624f
C71 top_c2.t2 VSUBS 3.7859f
C72 top_c2.n1 VSUBS 0.978608f
C73 top_c2.n2 VSUBS 0.909846f
C74 top_c0.t1 VSUBS 2.69371f
C75 top_c0.t0 VSUBS 2.48643f
C76 top_c0.n0 VSUBS 0.806119f
C77 top_c4.n0 VSUBS 0.068483f
C78 top_c4.n1 VSUBS 0.169865f
C79 top_c4.t13 VSUBS 1.93794f
C80 top_c4.n2 VSUBS 0.474158f
C81 top_c4.t1 VSUBS 1.07861f
C82 top_c4.n3 VSUBS 0.881063f
C83 top_c4.n4 VSUBS 0.41073f
C84 top_c4.n5 VSUBS 0.41073f
C85 top_c4.t11 VSUBS 1.07861f
C86 top_c4.n6 VSUBS 0.743495f
C87 top_c4.n7 VSUBS 0.150648f
C88 top_c4.t10 VSUBS 2.04439f
C89 top_c4.n8 VSUBS 0.210107f
C90 top_c4.t0 VSUBS 1.17567f
C91 top_c4.t9 VSUBS 1.85694f
C92 top_c4.n9 VSUBS 1.15519f
C93 top_c4.t7 VSUBS 1.07861f
C94 top_c4.n10 VSUBS 1.0908f
C95 top_c4.t8 VSUBS 1.07861f
C96 top_c4.n11 VSUBS 1.20383f
C97 top_c4.n12 VSUBS 0.251813f
C98 top_c4.t4 VSUBS 1.15435f
C99 top_c4.n13 VSUBS 1.1994f
C100 top_c4.n14 VSUBS 0.06994f
C101 top_c4.n15 VSUBS 0.06994f
C102 top_c4.t2 VSUBS 1.17567f
C103 top_c4.t14 VSUBS 1.85694f
C104 top_c4.n16 VSUBS 1.15519f
C105 top_c4.t12 VSUBS 1.07861f
C106 top_c4.n17 VSUBS 1.0908f
C107 top_c4.t3 VSUBS 1.07861f
C108 top_c4.n18 VSUBS 1.23178f
C109 top_c4.t6 VSUBS 2.09537f
C110 top_c4.n19 VSUBS 0.422503f
C111 top_c4.n20 VSUBS 0.152343f
C112 top_c4.t5 VSUBS 1.07861f
C113 top_c4.n21 VSUBS 0.76917f
C114 top_c4.n22 VSUBS 0.436457f
C115 top_c4.n23 VSUBS 0.436457f
C116 top_c4.t15 VSUBS 1.07861f
C117 top_c4.n24 VSUBS 0.500784f
C118 top_c4.n25 VSUBS 0.445419f
C119 top_c4.n26 VSUBS 0.088288f
C120 top_c4.n27 VSUBS 0.542953f
C121 top_c4.n28 VSUBS 0.623881f
C122 top_c3.t3 VSUBS 3.25884f
C123 top_c3.t0 VSUBS 3.03283f
C124 top_c3.n0 VSUBS 0.554743f
C125 top_c3.t1 VSUBS 2.95073f
C126 top_c3.n1 VSUBS 0.435391f
C127 top_c3.t7 VSUBS 3.03222f
C128 top_c3.n2 VSUBS 0.396406f
C129 top_c3.t4 VSUBS 3.004f
C130 top_c3.t6 VSUBS 3.09976f
C131 top_c3.n3 VSUBS 0.474775f
C132 top_c3.t2 VSUBS 2.95386f
C133 top_c3.n4 VSUBS 0.43584f
C134 top_c3.t5 VSUBS 3.21605f
C135 top_c3.n5 VSUBS 0.786601f
C136 top_c3.n6 VSUBS 0.632239f
C137 common_bottom.t51 VSUBS 1.10971f
C138 common_bottom.t28 VSUBS 1.18903f
C139 common_bottom.t52 VSUBS 1.19205f
C140 common_bottom.t38 VSUBS 1.1082f
C141 common_bottom.t5 VSUBS 1.18903f
C142 common_bottom.t44 VSUBS 1.18903f
C143 common_bottom.t7 VSUBS 1.19205f
C144 common_bottom.t58 VSUBS 1.18903f
C145 common_bottom.t16 VSUBS 1.19205f
C146 common_bottom.t57 VSUBS 1.18903f
C147 common_bottom.t49 VSUBS 1.19205f
C148 common_bottom.t59 VSUBS 1.19054f
C149 common_bottom.t0 VSUBS 1.19205f
C150 common_bottom.t26 VSUBS 1.10971f
C151 common_bottom.t12 VSUBS 1.10971f
C152 common_bottom.t47 VSUBS 1.18903f
C153 common_bottom.t25 VSUBS 1.1082f
C154 common_bottom.t39 VSUBS 1.03039f
C155 common_bottom.t61 VSUBS 1.18903f
C156 common_bottom.t27 VSUBS 1.18903f
C157 common_bottom.t13 VSUBS 1.18903f
C158 common_bottom.t41 VSUBS 1.10971f
C159 common_bottom.t10 VSUBS 1.10971f
C160 common_bottom.t43 VSUBS 1.10971f
C161 common_bottom.t9 VSUBS 1.10971f
C162 common_bottom.t23 VSUBS 1.10971f
C163 common_bottom.t11 VSUBS 1.18903f
C164 common_bottom.t62 VSUBS 1.19205f
C165 common_bottom.t15 VSUBS 1.10971f
C166 common_bottom.t37 VSUBS 1.10971f
C167 common_bottom.t18 VSUBS 1.18903f
C168 common_bottom.t36 VSUBS 1.19205f
C169 common_bottom.t20 VSUBS 1.19205f
C170 common_bottom.t3 VSUBS 1.18903f
C171 common_bottom.t46 VSUBS 1.18903f
C172 common_bottom.t8 VSUBS 1.19205f
C173 common_bottom.t54 VSUBS 1.10971f
C174 common_bottom.t50 VSUBS 1.02888f
C175 common_bottom.t2 VSUBS 1.11122f
C176 common_bottom.t42 VSUBS 1.1082f
C177 common_bottom.t30 VSUBS 1.1082f
C178 common_bottom.t40 VSUBS 1.11122f
C179 common_bottom.t33 VSUBS 1.11122f
C180 common_bottom.t19 VSUBS 1.1082f
C181 common_bottom.t35 VSUBS 1.02737f
C182 common_bottom.t22 VSUBS 1.11273f
C183 common_bottom.t24 VSUBS 1.1082f
C184 common_bottom.t53 VSUBS 1.19054f
C185 common_bottom.t1 VSUBS 1.19054f
C186 common_bottom.t45 VSUBS 1.19054f
C187 common_bottom.t21 VSUBS 1.19054f
C188 common_bottom.t55 VSUBS 1.19054f
C189 common_bottom.t63 VSUBS 1.19205f
C190 common_bottom.t31 VSUBS 1.19054f
C191 common_bottom.t48 VSUBS 1.18903f
C192 common_bottom.t60 VSUBS 1.19054f
C193 common_bottom.t14 VSUBS 1.19205f
C194 common_bottom.t29 VSUBS 1.19205f
C195 common_bottom.t4 VSUBS 1.19205f
C196 common_bottom.t32 VSUBS 1.19205f
C197 common_bottom.t17 VSUBS 1.11273f
C198 common_bottom.t34 VSUBS 1.10971f
C199 common_bottom.t56 VSUBS 1.1082f
C200 common_bottom.t6 VSUBS 1.10149f
C201 top_c5.n0 VSUBS 0.238348f
C202 top_c5.n1 VSUBS 0.265546f
C203 top_c5.n2 VSUBS 0.197079f
C204 top_c5.t21 VSUBS 0.668433f
C205 top_c5.n3 VSUBS 0.57654f
C206 top_c5.t3 VSUBS 0.668433f
C207 top_c5.n4 VSUBS 0.310344f
C208 top_c5.n5 VSUBS 0.217571f
C209 top_c5.t18 VSUBS 1.14806f
C210 top_c5.n6 VSUBS 0.332381f
C211 top_c5.t19 VSUBS 0.668433f
C212 top_c5.n7 VSUBS 0.310344f
C213 top_c5.n8 VSUBS 0.246374f
C214 top_c5.t9 VSUBS 0.668433f
C215 top_c5.n9 VSUBS 0.956132f
C216 top_c5.t31 VSUBS 0.668433f
C217 top_c5.n10 VSUBS 0.596691f
C218 top_c5.t7 VSUBS 0.668433f
C219 top_c5.n11 VSUBS 0.568189f
C220 top_c5.t5 VSUBS 1.21344f
C221 top_c5.n12 VSUBS 0.373736f
C222 top_c5.t22 VSUBS 0.668433f
C223 top_c5.n13 VSUBS 0.310344f
C224 top_c5.n14 VSUBS 0.276006f
C225 top_c5.t1 VSUBS 0.668433f
C226 top_c5.n15 VSUBS 0.717084f
C227 top_c5.t15 VSUBS 0.668433f
C228 top_c5.n16 VSUBS 0.717084f
C229 top_c5.n17 VSUBS 0.276833f
C230 top_c5.t17 VSUBS 0.668433f
C231 top_c5.n18 VSUBS 0.310344f
C232 top_c5.n19 VSUBS 0.264635f
C233 top_c5.t4 VSUBS 0.668433f
C234 top_c5.n20 VSUBS 0.310344f
C235 top_c5.n21 VSUBS 0.260893f
C236 top_c5.t20 VSUBS 0.668433f
C237 top_c5.n22 VSUBS 0.310344f
C238 top_c5.n23 VSUBS 0.189069f
C239 top_c5.t6 VSUBS 0.668433f
C240 top_c5.n24 VSUBS 0.473961f
C241 top_c5.n25 VSUBS 0.256817f
C242 top_c5.n26 VSUBS 0.263446f
C243 top_c5.n27 VSUBS 0.084591f
C244 top_c5.n28 VSUBS 0.072454f
C245 top_c5.n29 VSUBS 0.213794f
C246 top_c5.n30 VSUBS 0.265631f
C247 top_c5.t16 VSUBS 0.668433f
C248 top_c5.n31 VSUBS 0.315375f
C249 top_c5.t30 VSUBS 0.668433f
C250 top_c5.n32 VSUBS 0.439285f
C251 top_c5.n33 VSUBS 0.281344f
C252 top_c5.t28 VSUBS 0.668433f
C253 top_c5.n34 VSUBS 0.711294f
C254 top_c5.t8 VSUBS 0.668433f
C255 top_c5.n35 VSUBS 0.568189f
C256 top_c5.t2 VSUBS 1.27186f
C257 top_c5.n36 VSUBS 0.384211f
C258 top_c5.t24 VSUBS 0.668433f
C259 top_c5.n37 VSUBS 0.310344f
C260 top_c5.n38 VSUBS 0.276006f
C261 top_c5.t13 VSUBS 0.668433f
C262 top_c5.n39 VSUBS 0.717084f
C263 top_c5.t27 VSUBS 0.668433f
C264 top_c5.n40 VSUBS 0.717084f
C265 top_c5.n41 VSUBS 0.276006f
C266 top_c5.t14 VSUBS 0.668433f
C267 top_c5.n42 VSUBS 0.310344f
C268 top_c5.n43 VSUBS 0.268857f
C269 top_c5.n44 VSUBS 0.26096f
C270 top_c5.t0 VSUBS 0.668433f
C271 top_c5.n45 VSUBS 0.563401f
C272 top_c5.n46 VSUBS 0.08015f
C273 top_c5.n47 VSUBS 0.177877f
C274 top_c5.n48 VSUBS 0.218398f
C275 top_c5.t11 VSUBS 0.668433f
C276 top_c5.n49 VSUBS 0.69214f
C277 top_c5.t26 VSUBS 0.668433f
C278 top_c5.n50 VSUBS 0.310344f
C279 top_c5.n51 VSUBS 0.191012f
C280 top_c5.t10 VSUBS 0.728584f
C281 top_c5.t25 VSUBS 1.15077f
C282 top_c5.n52 VSUBS 0.715886f
C283 top_c5.t23 VSUBS 0.668433f
C284 top_c5.n53 VSUBS 0.665952f
C285 top_c5.n54 VSUBS 0.246374f
C286 top_c5.t12 VSUBS 0.668433f
C287 top_c5.n55 VSUBS 0.310344f
C288 top_c5.n56 VSUBS 0.246374f
C289 top_c5.t29 VSUBS 0.668433f
C290 top_c5.n57 VSUBS 0.645719f
C291 top_c5.n58 VSUBS 0.587047f
C292 top_c5.n59 VSUBS 0.48217f
.ends

