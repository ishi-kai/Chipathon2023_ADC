* NGSPICE file created from TOP.ext - technology: gf180mcuD

.subckt TOP VDD S R Q Qn GND
X0 GND.t56 Q.t30 Qn.t9 GND.t0 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X1 GND.t33 S.t0 Qn.t6 GND.t32 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X2 Qn.t15 Q.t31 GND.t55 GND.t30 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X3 Q.t5 Qn.t30 VDD.t19 VDD.t18 pfet_03v3 ad=0.728p pd=3.32u as=1.82p ps=6.9u w=2.8u l=0.28u
X4 VDD.t17 Qn.t31 Q.t9 VDD.t16 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X5 GND.t54 Q.t32 Qn.t14 GND.t4 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X6 GND.t42 R.t0 Q.t22 GND.t24 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X7 Q.t19 R.t1 GND.t39 GND.t20 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X8 VDD.t39 Q.t33 Qn.t27 VDD.t38 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X9 Q.t0 Qn.t32 VDD.t15 VDD.t14 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X10 VDD.t13 Qn.t33 Q.t3 VDD.t12 pfet_03v3 ad=1.82p pd=6.9u as=0.728p ps=3.32u w=2.8u l=0.28u
X11 Qn.t29 S.t1 GND.t59 GND.t49 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X12 GND.t25 Qn.t34 Q.t10 GND.t24 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X13 GND.t29 S.t2 Qn.t4 GND.t28 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X14 GND.t1 S.t3 Qn.t0 GND.t0 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X15 Q.t26 Qn.t35 GND.t23 GND.t22 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X16 Qn.t8 S.t4 GND.t45 GND.t44 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X17 Qn.t5 S.t5 GND.t31 GND.t30 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X18 Qn.t25 Q.t34 VDD.t37 VDD.t36 pfet_03v3 ad=0.728p pd=3.32u as=1.82p ps=6.9u w=2.8u l=0.28u
X19 VDD.t11 Qn.t36 Q.t2 VDD.t10 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X20 Q.t24 Qn.t37 GND.t21 GND.t20 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X21 Qn.t21 Q.t35 VDD.t35 VDD.t34 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X22 VDD.t33 Q.t36 Qn.t23 VDD.t32 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X23 GND.t19 Qn.t38 Q.t7 GND.t18 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X24 Q.t29 R.t2 GND.t58 GND.t16 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X25 Qn.t20 Q.t37 GND.t53 GND.t44 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X26 GND.t35 R.t3 Q.t14 GND.t12 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X27 GND.t34 R.t4 Q.t13 GND.t10 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X28 VDD.t9 Qn.t39 Q.t27 VDD.t8 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X29 Q.t23 R.t5 GND.t43 GND.t6 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X30 Q.t17 Qn.t40 VDD.t7 VDD.t6 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X31 GND.t52 Q.t38 Qn.t12 GND.t2 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X32 VDD.t31 Q.t39 Qn.t28 VDD.t30 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X33 Qn.t13 Q.t40 GND.t51 GND.t36 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X34 Qn.t17 Q.t41 GND.t50 GND.t49 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X35 GND.t3 S.t6 Qn.t1 GND.t2 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X36 GND.t48 Q.t42 Qn.t16 GND.t28 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X37 Qn.t7 S.t7 GND.t37 GND.t36 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X38 Q.t16 Qn.t41 VDD.t5 VDD.t4 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X39 Qn.t26 Q.t43 VDD.t29 VDD.t28 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X40 Q.t1 Qn.t42 GND.t17 GND.t16 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X41 Q.t11 Qn.t43 GND.t15 GND.t14 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X42 Q.t21 R.t6 GND.t41 GND.t22 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X43 VDD.t3 Qn.t44 Q.t15 VDD.t2 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X44 Q.t6 Qn.t45 VDD.t1 VDD.t0 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X45 GND.t38 R.t7 Q.t18 GND.t18 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X46 Qn.t22 Q.t44 VDD.t27 VDD.t26 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X47 VDD.t25 Q.t45 Qn.t24 VDD.t24 pfet_03v3 ad=1.82p pd=6.9u as=0.728p ps=3.32u w=2.8u l=0.28u
X48 GND.t13 Qn.t46 Q.t4 GND.t12 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X49 Q.t28 R.t8 GND.t57 GND.t14 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X50 GND.t11 Qn.t47 Q.t8 GND.t10 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X51 GND.t9 Qn.t48 Q.t12 GND.t8 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X52 GND.t40 R.t9 Q.t20 GND.t8 nfet_03v3 ad=1.708p pd=6.82u as=0.728p ps=3.32u w=2.8u l=0.28u
X53 Q.t25 Qn.t49 GND.t7 GND.t6 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X54 Qn.t19 Q.t46 GND.t47 GND.t26 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
X55 GND.t5 S.t8 Qn.t2 GND.t4 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X56 Qn.t18 Q.t47 VDD.t23 VDD.t22 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X57 GND.t46 Q.t48 Qn.t11 GND.t32 nfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X58 VDD.t21 Q.t49 Qn.t10 VDD.t20 pfet_03v3 ad=0.728p pd=3.32u as=0.728p ps=3.32u w=2.8u l=0.28u
X59 Qn.t3 S.t9 GND.t27 GND.t26 nfet_03v3 ad=0.728p pd=3.32u as=1.708p ps=6.82u w=2.8u l=0.28u
R0 Q.n0 Q.t45 55.9719
R1 Q.n1 Q.t34 55.9719
R2 Q.n2 Q.t33 55.9719
R3 Q.n3 Q.t43 55.9719
R4 Q.n4 Q.t39 55.9719
R5 Q.n5 Q.t35 55.9719
R6 Q.n6 Q.t49 55.9719
R7 Q.n7 Q.t44 55.9719
R8 Q.n8 Q.t36 55.9719
R9 Q.n9 Q.t47 55.9719
R10 Q.n1 Q.t46 55.9719
R11 Q.n2 Q.t48 55.9719
R12 Q.n3 Q.t37 55.9719
R13 Q.n4 Q.t30 55.9719
R14 Q.n5 Q.t31 55.9719
R15 Q.n6 Q.t38 55.9719
R16 Q.n7 Q.t40 55.9719
R17 Q.n8 Q.t32 55.9719
R18 Q.n9 Q.t41 55.9719
R19 Q.n0 Q.t42 55.9719
R20 Q.n35 Q.n21 7.35813
R21 Q.n33 Q.n22 7.35813
R22 Q.n31 Q.n23 7.35813
R23 Q.n29 Q.n24 7.35813
R24 Q.n27 Q.n25 7.35813
R25 Q.n13 Q.n11 5.94579
R26 Q.n35 Q.n34 5.90992
R27 Q.n33 Q.n32 5.90992
R28 Q.n31 Q.n30 5.90992
R29 Q.n29 Q.n28 5.90992
R30 Q.n27 Q.n26 5.90992
R31 Q.n20 Q.n10 5.71583
R32 Q.n19 Q.n18 5.69092
R33 Q.n17 Q.n16 5.69092
R34 Q.n15 Q.n14 5.69092
R35 Q.n13 Q.n12 5.69092
R36 Q.n18 Q.t27 0.6505
R37 Q.n18 Q.t5 0.6505
R38 Q.n16 Q.t9 0.6505
R39 Q.n16 Q.t16 0.6505
R40 Q.n14 Q.t15 0.6505
R41 Q.n14 Q.t17 0.6505
R42 Q.n12 Q.t2 0.6505
R43 Q.n12 Q.t0 0.6505
R44 Q.n11 Q.t3 0.6505
R45 Q.n11 Q.t6 0.6505
R46 Q.n34 Q.t4 0.5855
R47 Q.n34 Q.t26 0.5855
R48 Q.n21 Q.t14 0.5855
R49 Q.n21 Q.t21 0.5855
R50 Q.n32 Q.t10 0.5855
R51 Q.n32 Q.t1 0.5855
R52 Q.n22 Q.t22 0.5855
R53 Q.n22 Q.t29 0.5855
R54 Q.n30 Q.t7 0.5855
R55 Q.n30 Q.t11 0.5855
R56 Q.n23 Q.t18 0.5855
R57 Q.n23 Q.t28 0.5855
R58 Q.n28 Q.t8 0.5855
R59 Q.n28 Q.t25 0.5855
R60 Q.n24 Q.t13 0.5855
R61 Q.n24 Q.t23 0.5855
R62 Q.n26 Q.t12 0.5855
R63 Q.n26 Q.t24 0.5855
R64 Q.n25 Q.t20 0.5855
R65 Q.n25 Q.t19 0.5855
R66 Q.n20 Q.n19 0.39704
R67 Q Q.n35 0.271636
R68 Q.n15 Q.n13 0.255367
R69 Q.n17 Q.n15 0.255367
R70 Q.n19 Q.n17 0.255367
R71 Q.n29 Q.n27 0.223756
R72 Q.n31 Q.n29 0.223756
R73 Q.n33 Q.n31 0.223756
R74 Q.n35 Q.n33 0.223756
R75 Q.n9 Q.n8 0.0653649
R76 Q.n8 Q.n7 0.0653649
R77 Q.n7 Q.n6 0.0653649
R78 Q.n6 Q.n5 0.0653649
R79 Q.n5 Q.n4 0.0653649
R80 Q.n4 Q.n3 0.0653649
R81 Q.n3 Q.n2 0.0653649
R82 Q.n2 Q.n1 0.0653649
R83 Q.n10 Q.n0 0.0377911
R84 Q.n10 Q.n9 0.0288722
R85 Q Q.n20 0.0132703
R86 Qn.n9 Qn.t30 55.9719
R87 Qn.n8 Qn.t39 55.9719
R88 Qn.n7 Qn.t41 55.9719
R89 Qn.n6 Qn.t31 55.9719
R90 Qn.n5 Qn.t40 55.9719
R91 Qn.n4 Qn.t44 55.9719
R92 Qn.n3 Qn.t32 55.9719
R93 Qn.n2 Qn.t36 55.9719
R94 Qn.n1 Qn.t45 55.9719
R95 Qn.n0 Qn.t33 55.9719
R96 Qn.n9 Qn.t35 55.9719
R97 Qn.n8 Qn.t46 55.9719
R98 Qn.n7 Qn.t42 55.9719
R99 Qn.n6 Qn.t34 55.9719
R100 Qn.n5 Qn.t43 55.9719
R101 Qn.n4 Qn.t38 55.9719
R102 Qn.n3 Qn.t49 55.9719
R103 Qn.n2 Qn.t47 55.9719
R104 Qn.n1 Qn.t37 55.9719
R105 Qn.n0 Qn.t48 55.9719
R106 Qn.n27 Qn.n25 9.42441
R107 Qn.n29 Qn.n24 9.42441
R108 Qn.n31 Qn.n23 9.42441
R109 Qn.n33 Qn.n22 9.42441
R110 Qn.n35 Qn.n21 9.42441
R111 Qn.n27 Qn.n26 8.15873
R112 Qn.n29 Qn.n28 8.15873
R113 Qn.n31 Qn.n30 8.15873
R114 Qn.n33 Qn.n32 8.15873
R115 Qn.n35 Qn.n34 8.15873
R116 Qn.n13 Qn.n11 8.14399
R117 Qn.n13 Qn.n12 7.93973
R118 Qn.n15 Qn.n14 7.93973
R119 Qn.n17 Qn.n16 7.93973
R120 Qn.n19 Qn.n18 7.93973
R121 Qn.n20 Qn.n10 7.84476
R122 Qn.n11 Qn.t27 0.6505
R123 Qn.n11 Qn.t25 0.6505
R124 Qn.n12 Qn.t28 0.6505
R125 Qn.n12 Qn.t26 0.6505
R126 Qn.n14 Qn.t10 0.6505
R127 Qn.n14 Qn.t21 0.6505
R128 Qn.n16 Qn.t23 0.6505
R129 Qn.n16 Qn.t22 0.6505
R130 Qn.n18 Qn.t24 0.6505
R131 Qn.n18 Qn.t18 0.6505
R132 Qn.n26 Qn.t11 0.5855
R133 Qn.n26 Qn.t19 0.5855
R134 Qn.n25 Qn.t6 0.5855
R135 Qn.n25 Qn.t3 0.5855
R136 Qn.n28 Qn.t9 0.5855
R137 Qn.n28 Qn.t20 0.5855
R138 Qn.n24 Qn.t0 0.5855
R139 Qn.n24 Qn.t8 0.5855
R140 Qn.n30 Qn.t12 0.5855
R141 Qn.n30 Qn.t15 0.5855
R142 Qn.n23 Qn.t1 0.5855
R143 Qn.n23 Qn.t5 0.5855
R144 Qn.n32 Qn.t14 0.5855
R145 Qn.n32 Qn.t13 0.5855
R146 Qn.n22 Qn.t2 0.5855
R147 Qn.n22 Qn.t7 0.5855
R148 Qn.n34 Qn.t16 0.5855
R149 Qn.n34 Qn.t17 0.5855
R150 Qn.n21 Qn.t4 0.5855
R151 Qn.n21 Qn.t29 0.5855
R152 Qn Qn.n35 0.414192
R153 Qn.n20 Qn.n19 0.328301
R154 Qn.n35 Qn.n33 0.227272
R155 Qn.n33 Qn.n31 0.227272
R156 Qn.n31 Qn.n29 0.227272
R157 Qn.n29 Qn.n27 0.227272
R158 Qn.n19 Qn.n17 0.204755
R159 Qn.n17 Qn.n15 0.204755
R160 Qn.n15 Qn.n13 0.204755
R161 Qn.n1 Qn.n0 0.0653649
R162 Qn.n2 Qn.n1 0.0653649
R163 Qn.n3 Qn.n2 0.0653649
R164 Qn.n4 Qn.n3 0.0653649
R165 Qn.n5 Qn.n4 0.0653649
R166 Qn.n6 Qn.n5 0.0653649
R167 Qn.n7 Qn.n6 0.0653649
R168 Qn.n8 Qn.n7 0.0653649
R169 Qn.n10 Qn.n9 0.0357641
R170 Qn.n10 Qn.n8 0.0308992
R171 Qn Qn.n20 0.00161111
R172 GND.n29 GND.t8 25764.2
R173 GND.t26 GND.n29 25440.1
R174 GND.n29 GND.n17 8342.2
R175 GND.n28 GND.n17 575.247
R176 GND.n30 GND.n17 575.247
R177 GND.t22 GND.n28 365.005
R178 GND.n30 GND.t28 365.005
R179 GND.t8 GND.t20 233.603
R180 GND.t20 GND.t10 233.603
R181 GND.t10 GND.t6 233.603
R182 GND.t6 GND.t18 233.603
R183 GND.t18 GND.t14 233.603
R184 GND.t14 GND.t24 233.603
R185 GND.t24 GND.t16 233.603
R186 GND.t16 GND.t12 233.603
R187 GND.t12 GND.t22 233.603
R188 GND.t28 GND.t49 233.603
R189 GND.t49 GND.t4 233.603
R190 GND.t4 GND.t36 233.603
R191 GND.t36 GND.t2 233.603
R192 GND.t2 GND.t30 233.603
R193 GND.t30 GND.t0 233.603
R194 GND.t0 GND.t44 233.603
R195 GND.t44 GND.t32 233.603
R196 GND.t32 GND.t26 233.603
R197 GND.n18 GND.t23 9.84564
R198 GND.n6 GND.t9 9.83796
R199 GND.n18 GND.t41 9.05755
R200 GND.n6 GND.t40 9.05123
R201 GND.n5 GND.n3 8.94121
R202 GND.n2 GND.n0 8.94121
R203 GND.n24 GND.n22 8.94121
R204 GND.n21 GND.n19 8.94121
R205 GND.n5 GND.n4 8.15207
R206 GND.n2 GND.n1 8.15207
R207 GND.n24 GND.n23 8.15207
R208 GND.n21 GND.n20 8.15207
R209 GND.n40 GND.t47 7.60253
R210 GND.n16 GND.t48 7.60253
R211 GND.n16 GND.t29 6.81584
R212 GND.n40 GND.t27 6.81584
R213 GND.n15 GND.n13 6.70371
R214 GND.n12 GND.n10 6.70371
R215 GND.n36 GND.n34 6.70371
R216 GND.n39 GND.n37 6.70371
R217 GND.n15 GND.n14 5.91466
R218 GND.n12 GND.n11 5.91466
R219 GND.n36 GND.n35 5.91466
R220 GND.n39 GND.n38 5.91466
R221 GND.n28 GND.n27 5.59517
R222 GND.n31 GND.n30 4.56396
R223 GND.n41 GND.n40 1.07796
R224 GND.n7 GND.n6 0.991071
R225 GND.n31 GND.n16 0.899838
R226 GND.n32 GND.n15 0.898515
R227 GND.n33 GND.n12 0.898515
R228 GND.n42 GND.n36 0.898515
R229 GND.n41 GND.n39 0.898515
R230 GND.n7 GND.n5 0.862992
R231 GND.n8 GND.n2 0.862992
R232 GND.n25 GND.n24 0.862992
R233 GND.n26 GND.n21 0.862992
R234 GND.n27 GND.n18 0.862974
R235 GND GND.n9 0.66044
R236 GND.n4 GND.t39 0.5855
R237 GND.n4 GND.t34 0.5855
R238 GND.n3 GND.t21 0.5855
R239 GND.n3 GND.t11 0.5855
R240 GND.n1 GND.t43 0.5855
R241 GND.n1 GND.t38 0.5855
R242 GND.n0 GND.t7 0.5855
R243 GND.n0 GND.t19 0.5855
R244 GND.n23 GND.t57 0.5855
R245 GND.n23 GND.t42 0.5855
R246 GND.n22 GND.t15 0.5855
R247 GND.n22 GND.t25 0.5855
R248 GND.n20 GND.t58 0.5855
R249 GND.n20 GND.t35 0.5855
R250 GND.n19 GND.t17 0.5855
R251 GND.n19 GND.t13 0.5855
R252 GND.n14 GND.t59 0.5855
R253 GND.n14 GND.t5 0.5855
R254 GND.n13 GND.t50 0.5855
R255 GND.n13 GND.t54 0.5855
R256 GND.n11 GND.t37 0.5855
R257 GND.n11 GND.t3 0.5855
R258 GND.n10 GND.t51 0.5855
R259 GND.n10 GND.t52 0.5855
R260 GND.n35 GND.t31 0.5855
R261 GND.n35 GND.t1 0.5855
R262 GND.n34 GND.t55 0.5855
R263 GND.n34 GND.t56 0.5855
R264 GND.n38 GND.t45 0.5855
R265 GND.n38 GND.t33 0.5855
R266 GND.n37 GND.t53 0.5855
R267 GND.n37 GND.t46 0.5855
R268 GND GND.n43 0.503713
R269 GND.n32 GND.n31 0.143273
R270 GND.n33 GND.n32 0.131409
R271 GND.n42 GND.n41 0.131409
R272 GND.n27 GND.n26 0.12686
R273 GND.n8 GND.n7 0.1157
R274 GND.n26 GND.n25 0.1157
R275 GND.n43 GND.n42 0.0925455
R276 GND.n9 GND.n8 0.09086
R277 GND.n43 GND.n33 0.0393636
R278 GND.n25 GND.n9 0.02534
R279 S.n6 S.t9 56.1589
R280 S.n0 S.t2 56.1589
R281 S.n6 S.t0 55.9719
R282 S.n7 S.t4 55.9719
R283 S.n5 S.t3 55.9719
R284 S.n4 S.t5 55.9719
R285 S.n3 S.t6 55.9719
R286 S.n2 S.t7 55.9719
R287 S.n1 S.t8 55.9719
R288 S.n0 S.t1 55.9719
R289 S.n1 S.n0 0.187513
R290 S.n2 S.n1 0.187513
R291 S.n3 S.n2 0.187513
R292 S.n4 S.n3 0.187513
R293 S.n5 S.n4 0.187513
R294 S.n7 S.n6 0.187513
R295 S S.n5 0.106864
R296 S S.n7 0.0811494
R297 VDD.n6 VDD.t18 318.656
R298 VDD.n12 VDD.t24 316.43
R299 VDD.t0 VDD.t12 191.388
R300 VDD.t10 VDD.t0 191.388
R301 VDD.t14 VDD.t10 191.388
R302 VDD.t2 VDD.t14 191.388
R303 VDD.t6 VDD.t2 191.388
R304 VDD.t16 VDD.t6 191.388
R305 VDD.t4 VDD.t16 191.388
R306 VDD.t8 VDD.t4 191.388
R307 VDD.t18 VDD.t8 191.388
R308 VDD.t24 VDD.t22 191.388
R309 VDD.t22 VDD.t32 191.388
R310 VDD.t32 VDD.t26 191.388
R311 VDD.t26 VDD.t20 191.388
R312 VDD.t20 VDD.t34 191.388
R313 VDD.t34 VDD.t30 191.388
R314 VDD.t30 VDD.t28 191.388
R315 VDD.t28 VDD.t38 191.388
R316 VDD.t38 VDD.t36 191.388
R317 VDD.n2 VDD.t13 9.65475
R318 VDD.n6 VDD.t19 9.48844
R319 VDD.n7 VDD.n5 8.43844
R320 VDD.n8 VDD.n4 8.43844
R321 VDD.n3 VDD.n0 8.43844
R322 VDD.n2 VDD.n1 8.43844
R323 VDD.n17 VDD.t37 7.50384
R324 VDD.n12 VDD.t25 7.30419
R325 VDD.n17 VDD.n16 6.25419
R326 VDD.n18 VDD.n15 6.25419
R327 VDD.n14 VDD.n10 6.25419
R328 VDD.n13 VDD.n11 6.25419
R329 VDD VDD.n9 0.737162
R330 VDD.n5 VDD.t5 0.6505
R331 VDD.n5 VDD.t9 0.6505
R332 VDD.n4 VDD.t7 0.6505
R333 VDD.n4 VDD.t17 0.6505
R334 VDD.n0 VDD.t15 0.6505
R335 VDD.n0 VDD.t3 0.6505
R336 VDD.n1 VDD.t1 0.6505
R337 VDD.n1 VDD.t11 0.6505
R338 VDD.n16 VDD.t29 0.6505
R339 VDD.n16 VDD.t39 0.6505
R340 VDD.n15 VDD.t35 0.6505
R341 VDD.n15 VDD.t31 0.6505
R342 VDD.n10 VDD.t27 0.6505
R343 VDD.n10 VDD.t21 0.6505
R344 VDD.n11 VDD.t23 0.6505
R345 VDD.n11 VDD.t33 0.6505
R346 VDD VDD.n19 0.569824
R347 VDD.n7 VDD.n6 0.143273
R348 VDD.n13 VDD.n12 0.139447
R349 VDD.n3 VDD.n2 0.131409
R350 VDD.n8 VDD.n7 0.131409
R351 VDD.n14 VDD.n13 0.126816
R352 VDD.n18 VDD.n17 0.126816
R353 VDD.n19 VDD.n18 0.0983947
R354 VDD.n9 VDD.n3 0.0896818
R355 VDD.n9 VDD.n8 0.0422273
R356 VDD.n19 VDD.n14 0.0289211
R357 R.n4 R.t6 56.1655
R358 R.n0 R.t9 56.1655
R359 R.n7 R.t8 55.9719
R360 R.n6 R.t0 55.9719
R361 R.n5 R.t2 55.9719
R362 R.n4 R.t3 55.9719
R363 R.n3 R.t7 55.9719
R364 R.n2 R.t5 55.9719
R365 R.n1 R.t4 55.9719
R366 R.n0 R.t1 55.9719
R367 R.n5 R.n4 0.194062
R368 R.n6 R.n5 0.194062
R369 R.n7 R.n6 0.194062
R370 R.n1 R.n0 0.194062
R371 R.n2 R.n1 0.194062
R372 R.n3 R.n2 0.194062
R373 R R.n3 0.100979
R374 R R.n7 0.0935822
C0 Qn Q 3.31082f
C1 S VDD 0.013501f
C2 R Q 0.562407f
C3 Q VDD 5.65407f
C4 S Q 0.072343f
C5 R Qn 0.070425f
C6 Qn VDD 5.48142f
C7 R VDD 0.014082f
C8 S Qn 0.566319f
C9 R GND 2.73212f
C10 S GND 2.72481f
C11 Qn GND 12.066121f
C12 Q GND 12.538968f
C13 VDD GND 23.342003f
C14 VDD.t15 GND 0.021264f
C15 VDD.t3 GND 0.021264f
C16 VDD.n0 GND 0.11611f
C17 VDD.t1 GND 0.021264f
C18 VDD.t11 GND 0.021264f
C19 VDD.n1 GND 0.11611f
C20 VDD.t13 GND 0.166587f
C21 VDD.n2 GND 0.357459f
C22 VDD.n3 GND 0.172262f
C23 VDD.t7 GND 0.021264f
C24 VDD.t17 GND 0.021264f
C25 VDD.n4 GND 0.11611f
C26 VDD.t5 GND 0.021264f
C27 VDD.t9 GND 0.021264f
C28 VDD.n5 GND 0.11611f
C29 VDD.t19 GND 0.163795f
C30 VDD.t12 GND 0.459069f
C31 VDD.t0 GND 0.195349f
C32 VDD.t10 GND 0.195349f
C33 VDD.t14 GND 0.195349f
C34 VDD.t2 GND 0.195349f
C35 VDD.t6 GND 0.195349f
C36 VDD.t16 GND 0.195349f
C37 VDD.t4 GND 0.195349f
C38 VDD.t8 GND 0.195349f
C39 VDD.t18 GND 0.265946f
C40 VDD.n6 GND 0.620869f
C41 VDD.n7 GND 0.193307f
C42 VDD.n8 GND 0.153627f
C43 VDD.n9 GND 0.693672f
C44 VDD.t27 GND 0.021264f
C45 VDD.t21 GND 0.021264f
C46 VDD.n10 GND 0.102594f
C47 VDD.t23 GND 0.021264f
C48 VDD.t33 GND 0.021264f
C49 VDD.n11 GND 0.102594f
C50 VDD.t25 GND 0.147404f
C51 VDD.t36 GND 0.459069f
C52 VDD.t38 GND 0.195349f
C53 VDD.t28 GND 0.195349f
C54 VDD.t30 GND 0.195349f
C55 VDD.t34 GND 0.195349f
C56 VDD.t20 GND 0.195349f
C57 VDD.t26 GND 0.195349f
C58 VDD.t32 GND 0.195349f
C59 VDD.t22 GND 0.195349f
C60 VDD.t24 GND 0.263367f
C61 VDD.n12 GND 0.586909f
C62 VDD.n13 GND 0.181453f
C63 VDD.n14 GND 0.134836f
C64 VDD.t35 GND 0.021264f
C65 VDD.t31 GND 0.021264f
C66 VDD.n15 GND 0.102594f
C67 VDD.t29 GND 0.021264f
C68 VDD.t39 GND 0.021264f
C69 VDD.n16 GND 0.102594f
C70 VDD.t37 GND 0.150879f
C71 VDD.n17 GND 0.32623f
C72 VDD.n18 GND 0.164138f
C73 VDD.n19 GND 0.258997f
C74 Qn.t48 GND 0.051953f
C75 Qn.t33 GND 0.052152f
C76 Qn.n0 GND 0.104846f
C77 Qn.t37 GND 0.051953f
C78 Qn.t45 GND 0.052152f
C79 Qn.n1 GND 0.126076f
C80 Qn.t47 GND 0.051953f
C81 Qn.t36 GND 0.052152f
C82 Qn.n2 GND 0.126076f
C83 Qn.t49 GND 0.051953f
C84 Qn.t32 GND 0.052152f
C85 Qn.n3 GND 0.126076f
C86 Qn.t38 GND 0.051953f
C87 Qn.t44 GND 0.052152f
C88 Qn.n4 GND 0.126076f
C89 Qn.t43 GND 0.051953f
C90 Qn.t40 GND 0.052152f
C91 Qn.n5 GND 0.126076f
C92 Qn.t34 GND 0.051953f
C93 Qn.t31 GND 0.052152f
C94 Qn.n6 GND 0.126076f
C95 Qn.t42 GND 0.051953f
C96 Qn.t41 GND 0.052152f
C97 Qn.n7 GND 0.126076f
C98 Qn.t46 GND 0.051953f
C99 Qn.t39 GND 0.052152f
C100 Qn.n8 GND 0.115079f
C101 Qn.t35 GND 0.051953f
C102 Qn.t30 GND 0.052152f
C103 Qn.n9 GND 0.097942f
C104 Qn.n10 GND 0.077733f
C105 Qn.t27 GND 0.030691f
C106 Qn.t25 GND 0.030691f
C107 Qn.n11 GND 0.164422f
C108 Qn.t28 GND 0.030691f
C109 Qn.t26 GND 0.030691f
C110 Qn.n12 GND 0.161224f
C111 Qn.n13 GND 0.259499f
C112 Qn.t10 GND 0.030691f
C113 Qn.t21 GND 0.030691f
C114 Qn.n14 GND 0.161224f
C115 Qn.n15 GND 0.135212f
C116 Qn.t23 GND 0.030691f
C117 Qn.t22 GND 0.030691f
C118 Qn.n16 GND 0.161224f
C119 Qn.n17 GND 0.135212f
C120 Qn.t24 GND 0.030691f
C121 Qn.t18 GND 0.030691f
C122 Qn.n18 GND 0.161224f
C123 Qn.n19 GND 0.179245f
C124 Qn.n20 GND 0.323066f
C125 Qn.t4 GND 0.030691f
C126 Qn.t29 GND 0.030691f
C127 Qn.n21 GND 0.180762f
C128 Qn.t2 GND 0.030691f
C129 Qn.t7 GND 0.030691f
C130 Qn.n22 GND 0.180762f
C131 Qn.t1 GND 0.030691f
C132 Qn.t5 GND 0.030691f
C133 Qn.n23 GND 0.180762f
C134 Qn.t0 GND 0.030691f
C135 Qn.t8 GND 0.030691f
C136 Qn.n24 GND 0.180762f
C137 Qn.t6 GND 0.030691f
C138 Qn.t3 GND 0.030691f
C139 Qn.n25 GND 0.180762f
C140 Qn.t11 GND 0.030691f
C141 Qn.t19 GND 0.030691f
C142 Qn.n26 GND 0.158535f
C143 Qn.n27 GND 0.364671f
C144 Qn.t9 GND 0.030691f
C145 Qn.t20 GND 0.030691f
C146 Qn.n28 GND 0.158535f
C147 Qn.n29 GND 0.368151f
C148 Qn.t12 GND 0.030691f
C149 Qn.t15 GND 0.030691f
C150 Qn.n30 GND 0.158535f
C151 Qn.n31 GND 0.368151f
C152 Qn.t14 GND 0.030691f
C153 Qn.t13 GND 0.030691f
C154 Qn.n32 GND 0.158535f
C155 Qn.n33 GND 0.368151f
C156 Qn.t16 GND 0.030691f
C157 Qn.t17 GND 0.030691f
C158 Qn.n34 GND 0.158535f
C159 Qn.n35 GND 0.426811f
C160 Q.t42 GND 0.058973f
C161 Q.t45 GND 0.059198f
C162 Q.n0 GND 0.110814f
C163 Q.t41 GND 0.058973f
C164 Q.t32 GND 0.058973f
C165 Q.t40 GND 0.058973f
C166 Q.t38 GND 0.058973f
C167 Q.t31 GND 0.058973f
C168 Q.t30 GND 0.058973f
C169 Q.t37 GND 0.058973f
C170 Q.t48 GND 0.058973f
C171 Q.t46 GND 0.058973f
C172 Q.t34 GND 0.059198f
C173 Q.n1 GND 0.120802f
C174 Q.t33 GND 0.059198f
C175 Q.n2 GND 0.143112f
C176 Q.t43 GND 0.059198f
C177 Q.n3 GND 0.143112f
C178 Q.t39 GND 0.059198f
C179 Q.n4 GND 0.143112f
C180 Q.t35 GND 0.059198f
C181 Q.n5 GND 0.143112f
C182 Q.t49 GND 0.059198f
C183 Q.n6 GND 0.143112f
C184 Q.t44 GND 0.059198f
C185 Q.n7 GND 0.143112f
C186 Q.t36 GND 0.059198f
C187 Q.n8 GND 0.143112f
C188 Q.t47 GND 0.059198f
C189 Q.n9 GND 0.129819f
C190 Q.n10 GND 0.075577f
C191 Q.t3 GND 0.034838f
C192 Q.t6 GND 0.034838f
C193 Q.n11 GND 0.163629f
C194 Q.t2 GND 0.034838f
C195 Q.t0 GND 0.034838f
C196 Q.n12 GND 0.159308f
C197 Q.n13 GND 0.205112f
C198 Q.t15 GND 0.034838f
C199 Q.t17 GND 0.034838f
C200 Q.n14 GND 0.159308f
C201 Q.n15 GND 0.108637f
C202 Q.t9 GND 0.034838f
C203 Q.t16 GND 0.034838f
C204 Q.n16 GND 0.159308f
C205 Q.n17 GND 0.108637f
C206 Q.t27 GND 0.034838f
C207 Q.t5 GND 0.034838f
C208 Q.n18 GND 0.159308f
C209 Q.n19 GND 0.162941f
C210 Q.n20 GND 0.351105f
C211 Q.t14 GND 0.034838f
C212 Q.t21 GND 0.034838f
C213 Q.n21 GND 0.187432f
C214 Q.t22 GND 0.034838f
C215 Q.t29 GND 0.034838f
C216 Q.n22 GND 0.187432f
C217 Q.t18 GND 0.034838f
C218 Q.t28 GND 0.034838f
C219 Q.n23 GND 0.187432f
C220 Q.t13 GND 0.034838f
C221 Q.t23 GND 0.034838f
C222 Q.n24 GND 0.187432f
C223 Q.t20 GND 0.034838f
C224 Q.t19 GND 0.034838f
C225 Q.n25 GND 0.187432f
C226 Q.t12 GND 0.034838f
C227 Q.t24 GND 0.034838f
C228 Q.n26 GND 0.155972f
C229 Q.n27 GND 0.350142f
C230 Q.t8 GND 0.034838f
C231 Q.t25 GND 0.034838f
C232 Q.n28 GND 0.155972f
C233 Q.n29 GND 0.353538f
C234 Q.t7 GND 0.034838f
C235 Q.t11 GND 0.034838f
C236 Q.n30 GND 0.155972f
C237 Q.n31 GND 0.353538f
C238 Q.t10 GND 0.034838f
C239 Q.t1 GND 0.034838f
C240 Q.n32 GND 0.155972f
C241 Q.n33 GND 0.353538f
C242 Q.t4 GND 0.034838f
C243 Q.t26 GND 0.034838f
C244 Q.n34 GND 0.155972f
C245 Q.n35 GND 0.380023f
.ends

